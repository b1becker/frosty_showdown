library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity player1_rom is
	port(
		clk : in std_logic;
		x_cord : in unsigned(5 downto 0);
		y_cord : in unsigned(6 downto 0);
		rgb : out std_logic_vector(5 downto 0)
	);
end player1_rom;

architecture synth of player1_rom is
signal pxl : std_logic_vector(12 downto 0);
begin
	process(clk) begin
		if rising_edge(clk) then
			case pxl is	
            when "0000000000000" => rgb <= "100001";
            when "0000000000001" => rgb <= "100001";
            when "0000000000010" => rgb <= "100001";
            when "0000000000011" => rgb <= "100001";
            when "0000000000100" => rgb <= "100001";
            when "0000000000101" => rgb <= "100001";
            when "0000000000110" => rgb <= "100001";
            when "0000000000111" => rgb <= "100001";
            when "0000000001000" => rgb <= "100001";
            when "0000000001001" => rgb <= "100001";
            when "0000000001010" => rgb <= "100001";
            when "0000000001011" => rgb <= "100001";
            when "0000000001100" => rgb <= "100001";
            when "0000000001101" => rgb <= "000000";
            when "0000000001110" => rgb <= "000000";
            when "0000000001111" => rgb <= "000000";
            when "0000000010000" => rgb <= "000000";
            when "0000000010001" => rgb <= "000000";
            when "0000000010010" => rgb <= "000000";
            when "0000000010011" => rgb <= "000000";
            when "0000000010100" => rgb <= "000000";
            when "0000000010101" => rgb <= "000000";
            when "0000000010110" => rgb <= "000000";
            when "0000000010111" => rgb <= "000000";
            when "0000000011000" => rgb <= "000000";
            when "0000000011001" => rgb <= "000000";
            when "0000000011010" => rgb <= "000000";
            when "0000000011011" => rgb <= "000000";
            when "0000000011100" => rgb <= "000000";
            when "0000000011101" => rgb <= "100001";
            when "0000000011110" => rgb <= "100001";
            when "0000000011111" => rgb <= "100001";
            when "0000000100000" => rgb <= "100001";
            when "0000000100001" => rgb <= "100001";
            when "0000000100010" => rgb <= "100001";
            when "0000000100011" => rgb <= "100001";
            when "0000000100100" => rgb <= "100001";
            when "0000000100101" => rgb <= "100001";
            when "0000000100110" => rgb <= "100001";
            when "0000000100111" => rgb <= "100001";
            when "0000001000000" => rgb <= "100001";
            when "0000001000001" => rgb <= "100001";
            when "0000001000010" => rgb <= "100001";
            when "0000001000011" => rgb <= "100001";
            when "0000001000100" => rgb <= "100001";
            when "0000001000101" => rgb <= "100001";
            when "0000001000110" => rgb <= "100001";
            when "0000001000111" => rgb <= "100001";
            when "0000001001000" => rgb <= "100001";
            when "0000001001001" => rgb <= "100001";
            when "0000001001010" => rgb <= "100001";
            when "0000001001011" => rgb <= "100001";
            when "0000001001100" => rgb <= "100001";
            when "0000001001101" => rgb <= "000000";
            when "0000001001110" => rgb <= "000000";
            when "0000001001111" => rgb <= "000000";
            when "0000001010000" => rgb <= "000000";
            when "0000001010001" => rgb <= "000000";
            when "0000001010010" => rgb <= "000000";
            when "0000001010011" => rgb <= "000000";
            when "0000001010100" => rgb <= "000000";
            when "0000001010101" => rgb <= "000000";
            when "0000001010110" => rgb <= "000000";
            when "0000001010111" => rgb <= "000000";
            when "0000001011000" => rgb <= "000000";
            when "0000001011001" => rgb <= "000000";
            when "0000001011010" => rgb <= "000000";
            when "0000001011011" => rgb <= "000000";
            when "0000001011100" => rgb <= "000000";
            when "0000001011101" => rgb <= "100001";
            when "0000001011110" => rgb <= "100001";
            when "0000001011111" => rgb <= "100001";
            when "0000001100000" => rgb <= "100001";
            when "0000001100001" => rgb <= "100001";
            when "0000001100010" => rgb <= "100001";
            when "0000001100011" => rgb <= "100001";
            when "0000001100100" => rgb <= "100001";
            when "0000001100101" => rgb <= "100001";
            when "0000001100110" => rgb <= "100001";
            when "0000001100111" => rgb <= "100001";
            when "0000010000000" => rgb <= "100001";
            when "0000010000001" => rgb <= "100001";
            when "0000010000010" => rgb <= "100001";
            when "0000010000011" => rgb <= "100001";
            when "0000010000100" => rgb <= "100001";
            when "0000010000101" => rgb <= "100001";
            when "0000010000110" => rgb <= "100001";
            when "0000010000111" => rgb <= "100001";
            when "0000010001000" => rgb <= "100001";
            when "0000010001001" => rgb <= "100001";
            when "0000010001010" => rgb <= "100001";
            when "0000010001011" => rgb <= "100001";
            when "0000010001100" => rgb <= "100001";
            when "0000010001101" => rgb <= "000000";
            when "0000010001110" => rgb <= "000000";
            when "0000010001111" => rgb <= "000000";
            when "0000010010000" => rgb <= "000000";
            when "0000010010001" => rgb <= "000000";
            when "0000010010010" => rgb <= "000000";
            when "0000010010011" => rgb <= "000000";
            when "0000010010100" => rgb <= "000000";
            when "0000010010101" => rgb <= "000000";
            when "0000010010110" => rgb <= "000000";
            when "0000010010111" => rgb <= "000000";
            when "0000010011000" => rgb <= "000000";
            when "0000010011001" => rgb <= "000000";
            when "0000010011010" => rgb <= "000000";
            when "0000010011011" => rgb <= "000000";
            when "0000010011100" => rgb <= "000000";
            when "0000010011101" => rgb <= "100001";
            when "0000010011110" => rgb <= "100001";
            when "0000010011111" => rgb <= "100001";
            when "0000010100000" => rgb <= "100001";
            when "0000010100001" => rgb <= "100001";
            when "0000010100010" => rgb <= "100001";
            when "0000010100011" => rgb <= "100001";
            when "0000010100100" => rgb <= "100001";
            when "0000010100101" => rgb <= "100001";
            when "0000010100110" => rgb <= "100001";
            when "0000010100111" => rgb <= "100001";
            when "0000011000000" => rgb <= "100001";
            when "0000011000001" => rgb <= "100001";
            when "0000011000010" => rgb <= "100001";
            when "0000011000011" => rgb <= "100001";
            when "0000011000100" => rgb <= "100001";
            when "0000011000101" => rgb <= "100001";
            when "0000011000110" => rgb <= "100001";
            when "0000011000111" => rgb <= "100001";
            when "0000011001000" => rgb <= "100001";
            when "0000011001001" => rgb <= "100001";
            when "0000011001010" => rgb <= "100001";
            when "0000011001011" => rgb <= "100001";
            when "0000011001100" => rgb <= "100001";
            when "0000011001101" => rgb <= "000000";
            when "0000011001110" => rgb <= "000000";
            when "0000011001111" => rgb <= "000000";
            when "0000011010000" => rgb <= "000000";
            when "0000011010001" => rgb <= "000000";
            when "0000011010010" => rgb <= "000000";
            when "0000011010011" => rgb <= "000000";
            when "0000011010100" => rgb <= "000000";
            when "0000011010101" => rgb <= "000000";
            when "0000011010110" => rgb <= "000000";
            when "0000011010111" => rgb <= "000000";
            when "0000011011000" => rgb <= "000000";
            when "0000011011001" => rgb <= "000000";
            when "0000011011010" => rgb <= "000000";
            when "0000011011011" => rgb <= "000000";
            when "0000011011100" => rgb <= "000000";
            when "0000011011101" => rgb <= "100001";
            when "0000011011110" => rgb <= "100001";
            when "0000011011111" => rgb <= "100001";
            when "0000011100000" => rgb <= "100001";
            when "0000011100001" => rgb <= "100001";
            when "0000011100010" => rgb <= "100001";
            when "0000011100011" => rgb <= "100001";
            when "0000011100100" => rgb <= "100001";
            when "0000011100101" => rgb <= "100001";
            when "0000011100110" => rgb <= "100001";
            when "0000011100111" => rgb <= "100001";
            when "0000100000000" => rgb <= "100001";
            when "0000100000001" => rgb <= "100001";
            when "0000100000010" => rgb <= "100001";
            when "0000100000011" => rgb <= "100001";
            when "0000100000100" => rgb <= "100001";
            when "0000100000101" => rgb <= "100001";
            when "0000100000110" => rgb <= "100001";
            when "0000100000111" => rgb <= "100001";
            when "0000100001000" => rgb <= "100001";
            when "0000100001001" => rgb <= "100001";
            when "0000100001010" => rgb <= "100001";
            when "0000100001011" => rgb <= "100001";
            when "0000100001100" => rgb <= "100001";
            when "0000100001101" => rgb <= "000000";
            when "0000100001110" => rgb <= "000000";
            when "0000100001111" => rgb <= "000000";
            when "0000100010000" => rgb <= "000000";
            when "0000100010001" => rgb <= "000000";
            when "0000100010010" => rgb <= "000000";
            when "0000100010011" => rgb <= "000000";
            when "0000100010100" => rgb <= "000000";
            when "0000100010101" => rgb <= "000000";
            when "0000100010110" => rgb <= "000000";
            when "0000100010111" => rgb <= "000000";
            when "0000100011000" => rgb <= "000000";
            when "0000100011001" => rgb <= "000000";
            when "0000100011010" => rgb <= "000000";
            when "0000100011011" => rgb <= "000000";
            when "0000100011100" => rgb <= "000000";
            when "0000100011101" => rgb <= "100001";
            when "0000100011110" => rgb <= "100001";
            when "0000100011111" => rgb <= "100001";
            when "0000100100000" => rgb <= "100001";
            when "0000100100001" => rgb <= "100001";
            when "0000100100010" => rgb <= "100001";
            when "0000100100011" => rgb <= "100001";
            when "0000100100100" => rgb <= "100001";
            when "0000100100101" => rgb <= "100001";
            when "0000100100110" => rgb <= "100001";
            when "0000100100111" => rgb <= "100001";
            when "0000101000000" => rgb <= "100001";
            when "0000101000001" => rgb <= "100001";
            when "0000101000010" => rgb <= "100001";
            when "0000101000011" => rgb <= "100001";
            when "0000101000100" => rgb <= "100001";
            when "0000101000101" => rgb <= "100001";
            when "0000101000110" => rgb <= "100001";
            when "0000101000111" => rgb <= "100001";
            when "0000101001000" => rgb <= "100001";
            when "0000101001001" => rgb <= "100001";
            when "0000101001010" => rgb <= "100001";
            when "0000101001011" => rgb <= "100001";
            when "0000101001100" => rgb <= "100001";
            when "0000101001101" => rgb <= "000000";
            when "0000101001110" => rgb <= "000000";
            when "0000101001111" => rgb <= "000000";
            when "0000101010000" => rgb <= "000000";
            when "0000101010001" => rgb <= "000000";
            when "0000101010010" => rgb <= "000000";
            when "0000101010011" => rgb <= "000000";
            when "0000101010100" => rgb <= "000000";
            when "0000101010101" => rgb <= "000000";
            when "0000101010110" => rgb <= "000000";
            when "0000101010111" => rgb <= "000000";
            when "0000101011000" => rgb <= "000000";
            when "0000101011001" => rgb <= "000000";
            when "0000101011010" => rgb <= "000000";
            when "0000101011011" => rgb <= "000000";
            when "0000101011100" => rgb <= "000000";
            when "0000101011101" => rgb <= "100001";
            when "0000101011110" => rgb <= "100001";
            when "0000101011111" => rgb <= "100001";
            when "0000101100000" => rgb <= "100001";
            when "0000101100001" => rgb <= "100001";
            when "0000101100010" => rgb <= "100001";
            when "0000101100011" => rgb <= "100001";
            when "0000101100100" => rgb <= "100001";
            when "0000101100101" => rgb <= "100001";
            when "0000101100110" => rgb <= "100001";
            when "0000101100111" => rgb <= "100001";
            when "0000110000000" => rgb <= "100001";
            when "0000110000001" => rgb <= "100001";
            when "0000110000010" => rgb <= "100001";
            when "0000110000011" => rgb <= "100001";
            when "0000110000100" => rgb <= "100001";
            when "0000110000101" => rgb <= "100001";
            when "0000110000110" => rgb <= "100001";
            when "0000110000111" => rgb <= "100001";
            when "0000110001000" => rgb <= "100001";
            when "0000110001001" => rgb <= "100001";
            when "0000110001010" => rgb <= "100001";
            when "0000110001011" => rgb <= "100001";
            when "0000110001100" => rgb <= "100001";
            when "0000110001101" => rgb <= "000000";
            when "0000110001110" => rgb <= "000000";
            when "0000110001111" => rgb <= "000000";
            when "0000110010000" => rgb <= "000000";
            when "0000110010001" => rgb <= "000000";
            when "0000110010010" => rgb <= "000000";
            when "0000110010011" => rgb <= "000000";
            when "0000110010100" => rgb <= "000000";
            when "0000110010101" => rgb <= "000000";
            when "0000110010110" => rgb <= "000000";
            when "0000110010111" => rgb <= "000000";
            when "0000110011000" => rgb <= "000000";
            when "0000110011001" => rgb <= "000000";
            when "0000110011010" => rgb <= "000000";
            when "0000110011011" => rgb <= "000000";
            when "0000110011100" => rgb <= "000000";
            when "0000110011101" => rgb <= "100001";
            when "0000110011110" => rgb <= "100001";
            when "0000110011111" => rgb <= "100001";
            when "0000110100000" => rgb <= "100001";
            when "0000110100001" => rgb <= "100001";
            when "0000110100010" => rgb <= "100001";
            when "0000110100011" => rgb <= "100001";
            when "0000110100100" => rgb <= "100001";
            when "0000110100101" => rgb <= "100001";
            when "0000110100110" => rgb <= "100001";
            when "0000110100111" => rgb <= "100001";
            when "0000111000000" => rgb <= "100001";
            when "0000111000001" => rgb <= "100001";
            when "0000111000010" => rgb <= "100001";
            when "0000111000011" => rgb <= "100001";
            when "0000111000100" => rgb <= "100001";
            when "0000111000101" => rgb <= "100001";
            when "0000111000110" => rgb <= "100001";
            when "0000111000111" => rgb <= "100001";
            when "0000111001000" => rgb <= "100001";
            when "0000111001001" => rgb <= "100001";
            when "0000111001010" => rgb <= "100001";
            when "0000111001011" => rgb <= "100001";
            when "0000111001100" => rgb <= "100001";
            when "0000111001101" => rgb <= "000000";
            when "0000111001110" => rgb <= "000000";
            when "0000111001111" => rgb <= "000000";
            when "0000111010000" => rgb <= "000000";
            when "0000111010001" => rgb <= "000000";
            when "0000111010010" => rgb <= "000000";
            when "0000111010011" => rgb <= "000000";
            when "0000111010100" => rgb <= "000000";
            when "0000111010101" => rgb <= "000000";
            when "0000111010110" => rgb <= "000000";
            when "0000111010111" => rgb <= "000000";
            when "0000111011000" => rgb <= "000000";
            when "0000111011001" => rgb <= "000000";
            when "0000111011010" => rgb <= "000000";
            when "0000111011011" => rgb <= "000000";
            when "0000111011100" => rgb <= "000000";
            when "0000111011101" => rgb <= "100001";
            when "0000111011110" => rgb <= "100001";
            when "0000111011111" => rgb <= "100001";
            when "0000111100000" => rgb <= "100001";
            when "0000111100001" => rgb <= "100001";
            when "0000111100010" => rgb <= "100001";
            when "0000111100011" => rgb <= "100001";
            when "0000111100100" => rgb <= "100001";
            when "0000111100101" => rgb <= "100001";
            when "0000111100110" => rgb <= "100001";
            when "0000111100111" => rgb <= "100001";
            when "0001000000000" => rgb <= "100001";
            when "0001000000001" => rgb <= "100001";
            when "0001000000010" => rgb <= "100001";
            when "0001000000011" => rgb <= "100001";
            when "0001000000100" => rgb <= "100001";
            when "0001000000101" => rgb <= "100001";
            when "0001000000110" => rgb <= "100001";
            when "0001000000111" => rgb <= "100001";
            when "0001000001000" => rgb <= "100001";
            when "0001000001001" => rgb <= "100001";
            when "0001000001010" => rgb <= "100001";
            when "0001000001011" => rgb <= "100001";
            when "0001000001100" => rgb <= "100001";
            when "0001000001101" => rgb <= "000000";
            when "0001000001110" => rgb <= "000000";
            when "0001000001111" => rgb <= "000000";
            when "0001000010000" => rgb <= "000000";
            when "0001000010001" => rgb <= "000000";
            when "0001000010010" => rgb <= "000000";
            when "0001000010011" => rgb <= "000000";
            when "0001000010100" => rgb <= "000000";
            when "0001000010101" => rgb <= "000000";
            when "0001000010110" => rgb <= "000000";
            when "0001000010111" => rgb <= "000000";
            when "0001000011000" => rgb <= "000000";
            when "0001000011001" => rgb <= "000000";
            when "0001000011010" => rgb <= "000000";
            when "0001000011011" => rgb <= "000000";
            when "0001000011100" => rgb <= "000000";
            when "0001000011101" => rgb <= "100001";
            when "0001000011110" => rgb <= "100001";
            when "0001000011111" => rgb <= "100001";
            when "0001000100000" => rgb <= "100001";
            when "0001000100001" => rgb <= "100001";
            when "0001000100010" => rgb <= "100001";
            when "0001000100011" => rgb <= "100001";
            when "0001000100100" => rgb <= "100001";
            when "0001000100101" => rgb <= "100001";
            when "0001000100110" => rgb <= "100001";
            when "0001000100111" => rgb <= "100001";
            when "0001001000000" => rgb <= "100001";
            when "0001001000001" => rgb <= "100001";
            when "0001001000010" => rgb <= "100001";
            when "0001001000011" => rgb <= "100001";
            when "0001001000100" => rgb <= "100001";
            when "0001001000101" => rgb <= "100001";
            when "0001001000110" => rgb <= "100001";
            when "0001001000111" => rgb <= "100001";
            when "0001001001000" => rgb <= "100001";
            when "0001001001001" => rgb <= "100001";
            when "0001001001010" => rgb <= "100001";
            when "0001001001011" => rgb <= "100001";
            when "0001001001100" => rgb <= "100001";
            when "0001001001101" => rgb <= "000010";
            when "0001001001110" => rgb <= "000010";
            when "0001001001111" => rgb <= "000010";
            when "0001001010000" => rgb <= "000010";
            when "0001001010001" => rgb <= "000010";
            when "0001001010010" => rgb <= "000010";
            when "0001001010011" => rgb <= "000010";
            when "0001001010100" => rgb <= "000010";
            when "0001001010101" => rgb <= "000010";
            when "0001001010110" => rgb <= "000010";
            when "0001001010111" => rgb <= "000010";
            when "0001001011000" => rgb <= "000010";
            when "0001001011001" => rgb <= "000010";
            when "0001001011010" => rgb <= "000010";
            when "0001001011011" => rgb <= "000001";
            when "0001001011100" => rgb <= "000001";
            when "0001001011101" => rgb <= "100001";
            when "0001001011110" => rgb <= "100001";
            when "0001001011111" => rgb <= "100001";
            when "0001001100000" => rgb <= "100001";
            when "0001001100001" => rgb <= "100001";
            when "0001001100010" => rgb <= "100001";
            when "0001001100011" => rgb <= "100001";
            when "0001001100100" => rgb <= "100001";
            when "0001001100101" => rgb <= "100001";
            when "0001001100110" => rgb <= "100001";
            when "0001001100111" => rgb <= "100001";
            when "0001010000000" => rgb <= "100001";
            when "0001010000001" => rgb <= "100001";
            when "0001010000010" => rgb <= "100001";
            when "0001010000011" => rgb <= "100001";
            when "0001010000100" => rgb <= "100001";
            when "0001010000101" => rgb <= "100001";
            when "0001010000110" => rgb <= "100001";
            when "0001010000111" => rgb <= "100001";
            when "0001010001000" => rgb <= "100001";
            when "0001010001001" => rgb <= "100001";
            when "0001010001010" => rgb <= "100001";
            when "0001010001011" => rgb <= "100001";
            when "0001010001100" => rgb <= "100001";
            when "0001010001101" => rgb <= "000010";
            when "0001010001110" => rgb <= "000010";
            when "0001010001111" => rgb <= "000010";
            when "0001010010000" => rgb <= "000010";
            when "0001010010001" => rgb <= "000010";
            when "0001010010010" => rgb <= "000010";
            when "0001010010011" => rgb <= "000010";
            when "0001010010100" => rgb <= "000010";
            when "0001010010101" => rgb <= "000010";
            when "0001010010110" => rgb <= "000010";
            when "0001010010111" => rgb <= "000010";
            when "0001010011000" => rgb <= "000010";
            when "0001010011001" => rgb <= "000010";
            when "0001010011010" => rgb <= "000010";
            when "0001010011011" => rgb <= "000001";
            when "0001010011100" => rgb <= "000001";
            when "0001010011101" => rgb <= "100001";
            when "0001010011110" => rgb <= "100001";
            when "0001010011111" => rgb <= "100001";
            when "0001010100000" => rgb <= "100001";
            when "0001010100001" => rgb <= "100001";
            when "0001010100010" => rgb <= "100001";
            when "0001010100011" => rgb <= "100001";
            when "0001010100100" => rgb <= "100001";
            when "0001010100101" => rgb <= "100001";
            when "0001010100110" => rgb <= "100001";
            when "0001010100111" => rgb <= "100001";
            when "0001011000000" => rgb <= "100001";
            when "0001011000001" => rgb <= "100001";
            when "0001011000010" => rgb <= "100001";
            when "0001011000011" => rgb <= "100001";
            when "0001011000100" => rgb <= "100001";
            when "0001011000101" => rgb <= "100001";
            when "0001011000110" => rgb <= "100001";
            when "0001011000111" => rgb <= "100001";
            when "0001011001000" => rgb <= "100001";
            when "0001011001001" => rgb <= "100001";
            when "0001011001010" => rgb <= "100001";
            when "0001011001011" => rgb <= "100001";
            when "0001011001100" => rgb <= "100001";
            when "0001011001101" => rgb <= "000010";
            when "0001011001110" => rgb <= "000010";
            when "0001011001111" => rgb <= "000010";
            when "0001011010000" => rgb <= "000010";
            when "0001011010001" => rgb <= "000010";
            when "0001011010010" => rgb <= "000010";
            when "0001011010011" => rgb <= "000010";
            when "0001011010100" => rgb <= "000010";
            when "0001011010101" => rgb <= "000010";
            when "0001011010110" => rgb <= "000010";
            when "0001011010111" => rgb <= "000010";
            when "0001011011000" => rgb <= "000010";
            when "0001011011001" => rgb <= "000010";
            when "0001011011010" => rgb <= "000010";
            when "0001011011011" => rgb <= "000001";
            when "0001011011100" => rgb <= "000001";
            when "0001011011101" => rgb <= "100001";
            when "0001011011110" => rgb <= "100001";
            when "0001011011111" => rgb <= "100001";
            when "0001011100000" => rgb <= "100001";
            when "0001011100001" => rgb <= "100001";
            when "0001011100010" => rgb <= "100001";
            when "0001011100011" => rgb <= "100001";
            when "0001011100100" => rgb <= "100001";
            when "0001011100101" => rgb <= "100001";
            when "0001011100110" => rgb <= "100001";
            when "0001011100111" => rgb <= "100001";
            when "0001100000000" => rgb <= "100001";
            when "0001100000001" => rgb <= "100001";
            when "0001100000010" => rgb <= "100001";
            when "0001100000011" => rgb <= "100001";
            when "0001100000100" => rgb <= "100001";
            when "0001100000101" => rgb <= "100001";
            when "0001100000110" => rgb <= "100001";
            when "0001100000111" => rgb <= "100001";
            when "0001100001000" => rgb <= "100001";
            when "0001100001001" => rgb <= "100001";
            when "0001100001010" => rgb <= "100001";
            when "0001100001011" => rgb <= "100001";
            when "0001100001100" => rgb <= "100001";
            when "0001100001101" => rgb <= "000010";
            when "0001100001110" => rgb <= "000010";
            when "0001100001111" => rgb <= "000010";
            when "0001100010000" => rgb <= "000010";
            when "0001100010001" => rgb <= "000010";
            when "0001100010010" => rgb <= "000010";
            when "0001100010011" => rgb <= "000010";
            when "0001100010100" => rgb <= "000010";
            when "0001100010101" => rgb <= "000010";
            when "0001100010110" => rgb <= "000010";
            when "0001100010111" => rgb <= "000010";
            when "0001100011000" => rgb <= "000010";
            when "0001100011001" => rgb <= "000010";
            when "0001100011010" => rgb <= "000010";
            when "0001100011011" => rgb <= "000001";
            when "0001100011100" => rgb <= "000001";
            when "0001100011101" => rgb <= "100001";
            when "0001100011110" => rgb <= "100001";
            when "0001100011111" => rgb <= "100001";
            when "0001100100000" => rgb <= "100001";
            when "0001100100001" => rgb <= "100001";
            when "0001100100010" => rgb <= "100001";
            when "0001100100011" => rgb <= "100001";
            when "0001100100100" => rgb <= "100001";
            when "0001100100101" => rgb <= "100001";
            when "0001100100110" => rgb <= "100001";
            when "0001100100111" => rgb <= "100001";
            when "0001101000000" => rgb <= "100001";
            when "0001101000001" => rgb <= "100001";
            when "0001101000010" => rgb <= "100001";
            when "0001101000011" => rgb <= "100001";
            when "0001101000100" => rgb <= "100001";
            when "0001101000101" => rgb <= "100001";
            when "0001101000110" => rgb <= "100001";
            when "0001101000111" => rgb <= "100001";
            when "0001101001000" => rgb <= "100001";
            when "0001101001001" => rgb <= "100001";
            when "0001101001010" => rgb <= "100001";
            when "0001101001011" => rgb <= "100001";
            when "0001101001100" => rgb <= "000000";
            when "0001101001101" => rgb <= "000000";
            when "0001101001110" => rgb <= "000000";
            when "0001101001111" => rgb <= "000000";
            when "0001101010000" => rgb <= "000000";
            when "0001101010001" => rgb <= "000000";
            when "0001101010010" => rgb <= "000000";
            when "0001101010011" => rgb <= "000000";
            when "0001101010100" => rgb <= "000000";
            when "0001101010101" => rgb <= "000000";
            when "0001101010110" => rgb <= "000000";
            when "0001101010111" => rgb <= "000000";
            when "0001101011000" => rgb <= "000000";
            when "0001101011001" => rgb <= "000000";
            when "0001101011010" => rgb <= "000000";
            when "0001101011011" => rgb <= "000000";
            when "0001101011100" => rgb <= "000000";
            when "0001101011101" => rgb <= "000000";
            when "0001101011110" => rgb <= "100001";
            when "0001101011111" => rgb <= "100001";
            when "0001101100000" => rgb <= "100001";
            when "0001101100001" => rgb <= "100001";
            when "0001101100010" => rgb <= "100001";
            when "0001101100011" => rgb <= "100001";
            when "0001101100100" => rgb <= "100001";
            when "0001101100101" => rgb <= "100001";
            when "0001101100110" => rgb <= "100001";
            when "0001101100111" => rgb <= "100001";
            when "0001110000000" => rgb <= "100001";
            when "0001110000001" => rgb <= "100001";
            when "0001110000010" => rgb <= "100001";
            when "0001110000011" => rgb <= "100001";
            when "0001110000100" => rgb <= "100001";
            when "0001110000101" => rgb <= "100001";
            when "0001110000110" => rgb <= "100001";
            when "0001110000111" => rgb <= "100001";
            when "0001110001000" => rgb <= "100001";
            when "0001110001001" => rgb <= "100001";
            when "0001110001010" => rgb <= "100001";
            when "0001110001011" => rgb <= "100001";
            when "0001110001100" => rgb <= "000000";
            when "0001110001101" => rgb <= "000000";
            when "0001110001110" => rgb <= "000000";
            when "0001110001111" => rgb <= "000000";
            when "0001110010000" => rgb <= "000000";
            when "0001110010001" => rgb <= "000000";
            when "0001110010010" => rgb <= "000000";
            when "0001110010011" => rgb <= "000000";
            when "0001110010100" => rgb <= "000000";
            when "0001110010101" => rgb <= "000000";
            when "0001110010110" => rgb <= "000000";
            when "0001110010111" => rgb <= "000000";
            when "0001110011000" => rgb <= "000000";
            when "0001110011001" => rgb <= "000000";
            when "0001110011010" => rgb <= "000000";
            when "0001110011011" => rgb <= "000000";
            when "0001110011100" => rgb <= "000000";
            when "0001110011101" => rgb <= "000000";
            when "0001110011110" => rgb <= "100001";
            when "0001110011111" => rgb <= "100001";
            when "0001110100000" => rgb <= "100001";
            when "0001110100001" => rgb <= "100001";
            when "0001110100010" => rgb <= "100001";
            when "0001110100011" => rgb <= "100001";
            when "0001110100100" => rgb <= "100001";
            when "0001110100101" => rgb <= "100001";
            when "0001110100110" => rgb <= "100001";
            when "0001110100111" => rgb <= "100001";
            when "0001111000000" => rgb <= "100001";
            when "0001111000001" => rgb <= "100001";
            when "0001111000010" => rgb <= "100001";
            when "0001111000011" => rgb <= "100001";
            when "0001111000100" => rgb <= "100001";
            when "0001111000101" => rgb <= "100001";
            when "0001111000110" => rgb <= "100001";
            when "0001111000111" => rgb <= "100001";
            when "0001111001000" => rgb <= "100001";
            when "0001111001001" => rgb <= "100001";
            when "0001111001010" => rgb <= "100001";
            when "0001111001011" => rgb <= "100001";
            when "0001111001100" => rgb <= "000000";
            when "0001111001101" => rgb <= "000000";
            when "0001111001110" => rgb <= "000000";
            when "0001111001111" => rgb <= "000000";
            when "0001111010000" => rgb <= "000000";
            when "0001111010001" => rgb <= "000000";
            when "0001111010010" => rgb <= "000000";
            when "0001111010011" => rgb <= "000000";
            when "0001111010100" => rgb <= "000000";
            when "0001111010101" => rgb <= "000000";
            when "0001111010110" => rgb <= "000000";
            when "0001111010111" => rgb <= "000000";
            when "0001111011000" => rgb <= "000000";
            when "0001111011001" => rgb <= "000000";
            when "0001111011010" => rgb <= "000000";
            when "0001111011011" => rgb <= "000000";
            when "0001111011100" => rgb <= "000000";
            when "0001111011101" => rgb <= "000000";
            when "0001111011110" => rgb <= "100001";
            when "0001111011111" => rgb <= "100001";
            when "0001111100000" => rgb <= "100001";
            when "0001111100001" => rgb <= "100001";
            when "0001111100010" => rgb <= "100001";
            when "0001111100011" => rgb <= "100001";
            when "0001111100100" => rgb <= "100001";
            when "0001111100101" => rgb <= "100001";
            when "0001111100110" => rgb <= "100001";
            when "0001111100111" => rgb <= "100001";
            when "0010000000000" => rgb <= "100001";
            when "0010000000001" => rgb <= "100001";
            when "0010000000010" => rgb <= "100001";
            when "0010000000011" => rgb <= "100001";
            when "0010000000100" => rgb <= "100001";
            when "0010000000101" => rgb <= "100001";
            when "0010000000110" => rgb <= "100001";
            when "0010000000111" => rgb <= "100001";
            when "0010000001000" => rgb <= "100001";
            when "0010000001001" => rgb <= "100001";
            when "0010000001010" => rgb <= "100001";
            when "0010000001011" => rgb <= "100001";
            when "0010000001100" => rgb <= "000000";
            when "0010000001101" => rgb <= "000000";
            when "0010000001110" => rgb <= "000000";
            when "0010000001111" => rgb <= "000000";
            when "0010000010000" => rgb <= "000000";
            when "0010000010001" => rgb <= "000000";
            when "0010000010010" => rgb <= "000000";
            when "0010000010011" => rgb <= "000000";
            when "0010000010100" => rgb <= "000000";
            when "0010000010101" => rgb <= "000000";
            when "0010000010110" => rgb <= "000000";
            when "0010000010111" => rgb <= "000000";
            when "0010000011000" => rgb <= "000000";
            when "0010000011001" => rgb <= "000000";
            when "0010000011010" => rgb <= "000000";
            when "0010000011011" => rgb <= "000000";
            when "0010000011100" => rgb <= "000000";
            when "0010000011101" => rgb <= "000000";
            when "0010000011110" => rgb <= "100001";
            when "0010000011111" => rgb <= "100001";
            when "0010000100000" => rgb <= "100001";
            when "0010000100001" => rgb <= "100001";
            when "0010000100010" => rgb <= "100001";
            when "0010000100011" => rgb <= "100001";
            when "0010000100100" => rgb <= "100001";
            when "0010000100101" => rgb <= "100001";
            when "0010000100110" => rgb <= "100001";
            when "0010000100111" => rgb <= "100001";
            when "0010001000000" => rgb <= "100001";
            when "0010001000001" => rgb <= "100001";
            when "0010001000010" => rgb <= "100001";
            when "0010001000011" => rgb <= "100001";
            when "0010001000100" => rgb <= "100001";
            when "0010001000101" => rgb <= "100001";
            when "0010001000110" => rgb <= "100001";
            when "0010001000111" => rgb <= "100001";
            when "0010001001000" => rgb <= "000000";
            when "0010001001001" => rgb <= "000000";
            when "0010001001010" => rgb <= "000000";
            when "0010001001011" => rgb <= "000000";
            when "0010001001100" => rgb <= "000000";
            when "0010001001101" => rgb <= "000000";
            when "0010001001110" => rgb <= "000000";
            when "0010001001111" => rgb <= "000000";
            when "0010001010000" => rgb <= "000000";
            when "0010001010001" => rgb <= "000000";
            when "0010001010010" => rgb <= "000000";
            when "0010001010011" => rgb <= "000000";
            when "0010001010100" => rgb <= "000000";
            when "0010001010101" => rgb <= "000000";
            when "0010001010110" => rgb <= "000000";
            when "0010001010111" => rgb <= "000000";
            when "0010001011000" => rgb <= "000000";
            when "0010001011001" => rgb <= "000000";
            when "0010001011010" => rgb <= "000000";
            when "0010001011011" => rgb <= "000000";
            when "0010001011100" => rgb <= "000000";
            when "0010001011101" => rgb <= "000000";
            when "0010001011110" => rgb <= "000000";
            when "0010001011111" => rgb <= "000000";
            when "0010001100000" => rgb <= "000000";
            when "0010001100001" => rgb <= "000000";
            when "0010001100010" => rgb <= "100001";
            when "0010001100011" => rgb <= "100001";
            when "0010001100100" => rgb <= "100001";
            when "0010001100101" => rgb <= "100001";
            when "0010001100110" => rgb <= "100001";
            when "0010001100111" => rgb <= "100001";
            when "0010010000000" => rgb <= "100001";
            when "0010010000001" => rgb <= "100001";
            when "0010010000010" => rgb <= "100001";
            when "0010010000011" => rgb <= "100001";
            when "0010010000100" => rgb <= "100001";
            when "0010010000101" => rgb <= "100001";
            when "0010010000110" => rgb <= "100001";
            when "0010010000111" => rgb <= "100001";
            when "0010010001000" => rgb <= "000000";
            when "0010010001001" => rgb <= "000000";
            when "0010010001010" => rgb <= "000000";
            when "0010010001011" => rgb <= "000000";
            when "0010010001100" => rgb <= "000000";
            when "0010010001101" => rgb <= "000000";
            when "0010010001110" => rgb <= "000000";
            when "0010010001111" => rgb <= "000000";
            when "0010010010000" => rgb <= "000000";
            when "0010010010001" => rgb <= "000000";
            when "0010010010010" => rgb <= "000000";
            when "0010010010011" => rgb <= "000000";
            when "0010010010100" => rgb <= "000000";
            when "0010010010101" => rgb <= "000000";
            when "0010010010110" => rgb <= "000000";
            when "0010010010111" => rgb <= "000000";
            when "0010010011000" => rgb <= "000000";
            when "0010010011001" => rgb <= "000000";
            when "0010010011010" => rgb <= "000000";
            when "0010010011011" => rgb <= "000000";
            when "0010010011100" => rgb <= "000000";
            when "0010010011101" => rgb <= "000000";
            when "0010010011110" => rgb <= "000000";
            when "0010010011111" => rgb <= "000000";
            when "0010010100000" => rgb <= "000000";
            when "0010010100001" => rgb <= "000000";
            when "0010010100010" => rgb <= "100001";
            when "0010010100011" => rgb <= "100001";
            when "0010010100100" => rgb <= "100001";
            when "0010010100101" => rgb <= "100001";
            when "0010010100110" => rgb <= "100001";
            when "0010010100111" => rgb <= "100001";
            when "0010011000000" => rgb <= "100001";
            when "0010011000001" => rgb <= "100001";
            when "0010011000010" => rgb <= "100001";
            when "0010011000011" => rgb <= "100001";
            when "0010011000100" => rgb <= "100001";
            when "0010011000101" => rgb <= "100001";
            when "0010011000110" => rgb <= "100001";
            when "0010011000111" => rgb <= "100001";
            when "0010011001000" => rgb <= "100001";
            when "0010011001001" => rgb <= "100001";
            when "0010011001010" => rgb <= "100001";
            when "0010011001011" => rgb <= "010101";
            when "0010011001100" => rgb <= "101010";
            when "0010011001101" => rgb <= "101010";
            when "0010011001110" => rgb <= "101010";
            when "0010011001111" => rgb <= "101010";
            when "0010011010000" => rgb <= "101010";
            when "0010011010001" => rgb <= "111111";
            when "0010011010010" => rgb <= "111111";
            when "0010011010011" => rgb <= "111111";
            when "0010011010100" => rgb <= "111111";
            when "0010011010101" => rgb <= "111111";
            when "0010011010110" => rgb <= "111111";
            when "0010011010111" => rgb <= "111111";
            when "0010011011000" => rgb <= "111111";
            when "0010011011001" => rgb <= "111111";
            when "0010011011010" => rgb <= "111111";
            when "0010011011011" => rgb <= "111111";
            when "0010011011100" => rgb <= "111111";
            when "0010011011101" => rgb <= "010101";
            when "0010011011110" => rgb <= "100001";
            when "0010011011111" => rgb <= "100001";
            when "0010011100000" => rgb <= "100001";
            when "0010011100001" => rgb <= "100001";
            when "0010011100010" => rgb <= "100001";
            when "0010011100011" => rgb <= "100001";
            when "0010011100100" => rgb <= "100001";
            when "0010011100101" => rgb <= "100001";
            when "0010011100110" => rgb <= "100001";
            when "0010011100111" => rgb <= "100001";
            when "0010100000000" => rgb <= "100001";
            when "0010100000001" => rgb <= "100001";
            when "0010100000010" => rgb <= "100001";
            when "0010100000011" => rgb <= "100001";
            when "0010100000100" => rgb <= "100001";
            when "0010100000101" => rgb <= "100001";
            when "0010100000110" => rgb <= "100001";
            when "0010100000111" => rgb <= "100001";
            when "0010100001000" => rgb <= "100001";
            when "0010100001001" => rgb <= "100001";
            when "0010100001010" => rgb <= "100001";
            when "0010100001011" => rgb <= "010101";
            when "0010100001100" => rgb <= "101010";
            when "0010100001101" => rgb <= "101010";
            when "0010100001110" => rgb <= "101010";
            when "0010100001111" => rgb <= "101010";
            when "0010100010000" => rgb <= "101010";
            when "0010100010001" => rgb <= "111111";
            when "0010100010010" => rgb <= "111111";
            when "0010100010011" => rgb <= "111111";
            when "0010100010100" => rgb <= "111111";
            when "0010100010101" => rgb <= "111111";
            when "0010100010110" => rgb <= "111111";
            when "0010100010111" => rgb <= "111111";
            when "0010100011000" => rgb <= "111111";
            when "0010100011001" => rgb <= "111111";
            when "0010100011010" => rgb <= "111111";
            when "0010100011011" => rgb <= "111111";
            when "0010100011100" => rgb <= "111111";
            when "0010100011101" => rgb <= "010101";
            when "0010100011110" => rgb <= "100001";
            when "0010100011111" => rgb <= "100001";
            when "0010100100000" => rgb <= "100001";
            when "0010100100001" => rgb <= "100001";
            when "0010100100010" => rgb <= "100001";
            when "0010100100011" => rgb <= "100001";
            when "0010100100100" => rgb <= "100001";
            when "0010100100101" => rgb <= "100001";
            when "0010100100110" => rgb <= "100001";
            when "0010100100111" => rgb <= "100001";
            when "0010101000000" => rgb <= "100001";
            when "0010101000001" => rgb <= "100001";
            when "0010101000010" => rgb <= "100001";
            when "0010101000011" => rgb <= "100001";
            when "0010101000100" => rgb <= "100001";
            when "0010101000101" => rgb <= "100001";
            when "0010101000110" => rgb <= "100001";
            when "0010101000111" => rgb <= "100001";
            when "0010101001000" => rgb <= "100001";
            when "0010101001001" => rgb <= "100001";
            when "0010101001010" => rgb <= "010101";
            when "0010101001011" => rgb <= "101010";
            when "0010101001100" => rgb <= "101010";
            when "0010101001101" => rgb <= "101010";
            when "0010101001110" => rgb <= "111111";
            when "0010101001111" => rgb <= "111111";
            when "0010101010000" => rgb <= "111111";
            when "0010101010001" => rgb <= "111111";
            when "0010101010010" => rgb <= "111111";
            when "0010101010011" => rgb <= "111111";
            when "0010101010100" => rgb <= "111111";
            when "0010101010101" => rgb <= "111111";
            when "0010101010110" => rgb <= "111111";
            when "0010101010111" => rgb <= "111111";
            when "0010101011000" => rgb <= "111111";
            when "0010101011001" => rgb <= "111111";
            when "0010101011010" => rgb <= "111111";
            when "0010101011011" => rgb <= "111111";
            when "0010101011100" => rgb <= "111111";
            when "0010101011101" => rgb <= "111111";
            when "0010101011110" => rgb <= "010101";
            when "0010101011111" => rgb <= "100001";
            when "0010101100000" => rgb <= "100001";
            when "0010101100001" => rgb <= "100001";
            when "0010101100010" => rgb <= "100001";
            when "0010101100011" => rgb <= "100001";
            when "0010101100100" => rgb <= "100001";
            when "0010101100101" => rgb <= "100001";
            when "0010101100110" => rgb <= "100001";
            when "0010101100111" => rgb <= "100001";
            when "0010110000000" => rgb <= "100001";
            when "0010110000001" => rgb <= "100001";
            when "0010110000010" => rgb <= "100001";
            when "0010110000011" => rgb <= "100001";
            when "0010110000100" => rgb <= "100001";
            when "0010110000101" => rgb <= "100001";
            when "0010110000110" => rgb <= "100001";
            when "0010110000111" => rgb <= "100001";
            when "0010110001000" => rgb <= "100001";
            when "0010110001001" => rgb <= "010101";
            when "0010110001010" => rgb <= "101010";
            when "0010110001011" => rgb <= "101010";
            when "0010110001100" => rgb <= "111111";
            when "0010110001101" => rgb <= "111111";
            when "0010110001110" => rgb <= "111111";
            when "0010110001111" => rgb <= "111111";
            when "0010110010000" => rgb <= "111111";
            when "0010110010001" => rgb <= "111111";
            when "0010110010010" => rgb <= "111111";
            when "0010110010011" => rgb <= "111111";
            when "0010110010100" => rgb <= "111111";
            when "0010110010101" => rgb <= "111111";
            when "0010110010110" => rgb <= "111111";
            when "0010110010111" => rgb <= "111111";
            when "0010110011000" => rgb <= "111111";
            when "0010110011001" => rgb <= "111111";
            when "0010110011010" => rgb <= "111111";
            when "0010110011011" => rgb <= "111111";
            when "0010110011100" => rgb <= "111111";
            when "0010110011101" => rgb <= "111111";
            when "0010110011110" => rgb <= "111111";
            when "0010110011111" => rgb <= "010101";
            when "0010110100000" => rgb <= "100001";
            when "0010110100001" => rgb <= "100001";
            when "0010110100010" => rgb <= "100001";
            when "0010110100011" => rgb <= "100001";
            when "0010110100100" => rgb <= "100001";
            when "0010110100101" => rgb <= "100001";
            when "0010110100110" => rgb <= "100001";
            when "0010110100111" => rgb <= "100001";
            when "0010111000000" => rgb <= "100001";
            when "0010111000001" => rgb <= "100001";
            when "0010111000010" => rgb <= "100001";
            when "0010111000011" => rgb <= "100001";
            when "0010111000100" => rgb <= "100001";
            when "0010111000101" => rgb <= "100001";
            when "0010111000110" => rgb <= "100001";
            when "0010111000111" => rgb <= "100001";
            when "0010111001000" => rgb <= "010101";
            when "0010111001001" => rgb <= "101010";
            when "0010111001010" => rgb <= "101010";
            when "0010111001011" => rgb <= "111111";
            when "0010111001100" => rgb <= "111111";
            when "0010111001101" => rgb <= "111111";
            when "0010111001110" => rgb <= "111111";
            when "0010111001111" => rgb <= "111111";
            when "0010111010000" => rgb <= "111111";
            when "0010111010001" => rgb <= "111111";
            when "0010111010010" => rgb <= "111111";
            when "0010111010011" => rgb <= "111111";
            when "0010111010100" => rgb <= "111111";
            when "0010111010101" => rgb <= "111111";
            when "0010111010110" => rgb <= "111111";
            when "0010111010111" => rgb <= "111111";
            when "0010111011000" => rgb <= "111111";
            when "0010111011001" => rgb <= "111111";
            when "0010111011010" => rgb <= "111111";
            when "0010111011011" => rgb <= "111111";
            when "0010111011100" => rgb <= "111111";
            when "0010111011101" => rgb <= "111111";
            when "0010111011110" => rgb <= "111111";
            when "0010111011111" => rgb <= "111111";
            when "0010111100000" => rgb <= "010101";
            when "0010111100001" => rgb <= "100001";
            when "0010111100010" => rgb <= "100001";
            when "0010111100011" => rgb <= "100001";
            when "0010111100100" => rgb <= "100001";
            when "0010111100101" => rgb <= "100001";
            when "0010111100110" => rgb <= "100001";
            when "0010111100111" => rgb <= "100001";
            when "0011000000000" => rgb <= "100001";
            when "0011000000001" => rgb <= "100001";
            when "0011000000010" => rgb <= "100001";
            when "0011000000011" => rgb <= "100001";
            when "0011000000100" => rgb <= "100001";
            when "0011000000101" => rgb <= "100001";
            when "0011000000110" => rgb <= "100001";
            when "0011000000111" => rgb <= "100001";
            when "0011000001000" => rgb <= "010101";
            when "0011000001001" => rgb <= "101010";
            when "0011000001010" => rgb <= "101010";
            when "0011000001011" => rgb <= "111111";
            when "0011000001100" => rgb <= "111111";
            when "0011000001101" => rgb <= "111111";
            when "0011000001110" => rgb <= "111111";
            when "0011000001111" => rgb <= "111111";
            when "0011000010000" => rgb <= "111111";
            when "0011000010001" => rgb <= "111111";
            when "0011000010010" => rgb <= "111111";
            when "0011000010011" => rgb <= "111111";
            when "0011000010100" => rgb <= "111111";
            when "0011000010101" => rgb <= "111111";
            when "0011000010110" => rgb <= "111111";
            when "0011000010111" => rgb <= "111111";
            when "0011000011000" => rgb <= "111111";
            when "0011000011001" => rgb <= "111111";
            when "0011000011010" => rgb <= "111111";
            when "0011000011011" => rgb <= "111111";
            when "0011000011100" => rgb <= "111111";
            when "0011000011101" => rgb <= "111111";
            when "0011000011110" => rgb <= "111111";
            when "0011000011111" => rgb <= "111111";
            when "0011000100000" => rgb <= "010101";
            when "0011000100001" => rgb <= "100001";
            when "0011000100010" => rgb <= "100001";
            when "0011000100011" => rgb <= "100001";
            when "0011000100100" => rgb <= "100001";
            when "0011000100101" => rgb <= "100001";
            when "0011000100110" => rgb <= "100001";
            when "0011000100111" => rgb <= "100001";
            when "0011001000000" => rgb <= "100001";
            when "0011001000001" => rgb <= "100001";
            when "0011001000010" => rgb <= "100001";
            when "0011001000011" => rgb <= "100001";
            when "0011001000100" => rgb <= "100001";
            when "0011001000101" => rgb <= "100001";
            when "0011001000110" => rgb <= "100001";
            when "0011001000111" => rgb <= "100001";
            when "0011001001000" => rgb <= "010101";
            when "0011001001001" => rgb <= "101010";
            when "0011001001010" => rgb <= "101010";
            when "0011001001011" => rgb <= "111111";
            when "0011001001100" => rgb <= "111111";
            when "0011001001101" => rgb <= "111111";
            when "0011001001110" => rgb <= "111111";
            when "0011001001111" => rgb <= "111111";
            when "0011001010000" => rgb <= "111111";
            when "0011001010001" => rgb <= "111111";
            when "0011001010010" => rgb <= "111111";
            when "0011001010011" => rgb <= "111111";
            when "0011001010100" => rgb <= "111111";
            when "0011001010101" => rgb <= "111111";
            when "0011001010110" => rgb <= "111111";
            when "0011001010111" => rgb <= "111111";
            when "0011001011000" => rgb <= "111111";
            when "0011001011001" => rgb <= "111111";
            when "0011001011010" => rgb <= "111111";
            when "0011001011011" => rgb <= "111111";
            when "0011001011100" => rgb <= "111111";
            when "0011001011101" => rgb <= "111111";
            when "0011001011110" => rgb <= "111111";
            when "0011001011111" => rgb <= "111111";
            when "0011001100000" => rgb <= "010101";
            when "0011001100001" => rgb <= "100001";
            when "0011001100010" => rgb <= "100001";
            when "0011001100011" => rgb <= "100001";
            when "0011001100100" => rgb <= "100001";
            when "0011001100101" => rgb <= "100001";
            when "0011001100110" => rgb <= "100001";
            when "0011001100111" => rgb <= "100001";
            when "0011010000000" => rgb <= "100001";
            when "0011010000001" => rgb <= "100001";
            when "0011010000010" => rgb <= "100001";
            when "0011010000011" => rgb <= "100001";
            when "0011010000100" => rgb <= "100001";
            when "0011010000101" => rgb <= "100001";
            when "0011010000110" => rgb <= "100001";
            when "0011010000111" => rgb <= "010101";
            when "0011010001000" => rgb <= "101010";
            when "0011010001001" => rgb <= "101010";
            when "0011010001010" => rgb <= "111111";
            when "0011010001011" => rgb <= "111111";
            when "0011010001100" => rgb <= "111111";
            when "0011010001101" => rgb <= "111111";
            when "0011010001110" => rgb <= "111111";
            when "0011010001111" => rgb <= "111111";
            when "0011010010000" => rgb <= "111111";
            when "0011010010001" => rgb <= "111111";
            when "0011010010010" => rgb <= "111111";
            when "0011010010011" => rgb <= "111111";
            when "0011010010100" => rgb <= "111111";
            when "0011010010101" => rgb <= "111111";
            when "0011010010110" => rgb <= "111111";
            when "0011010010111" => rgb <= "111111";
            when "0011010011000" => rgb <= "111111";
            when "0011010011001" => rgb <= "111111";
            when "0011010011010" => rgb <= "111111";
            when "0011010011011" => rgb <= "111111";
            when "0011010011100" => rgb <= "111111";
            when "0011010011101" => rgb <= "111111";
            when "0011010011110" => rgb <= "111111";
            when "0011010011111" => rgb <= "111111";
            when "0011010100000" => rgb <= "111111";
            when "0011010100001" => rgb <= "010101";
            when "0011010100010" => rgb <= "100001";
            when "0011010100011" => rgb <= "100001";
            when "0011010100100" => rgb <= "100001";
            when "0011010100101" => rgb <= "100001";
            when "0011010100110" => rgb <= "100001";
            when "0011010100111" => rgb <= "100001";
            when "0011011000000" => rgb <= "100001";
            when "0011011000001" => rgb <= "100001";
            when "0011011000010" => rgb <= "100001";
            when "0011011000011" => rgb <= "100001";
            when "0011011000100" => rgb <= "100001";
            when "0011011000101" => rgb <= "100001";
            when "0011011000110" => rgb <= "100001";
            when "0011011000111" => rgb <= "010101";
            when "0011011001000" => rgb <= "101010";
            when "0011011001001" => rgb <= "101010";
            when "0011011001010" => rgb <= "111111";
            when "0011011001011" => rgb <= "111111";
            when "0011011001100" => rgb <= "111111";
            when "0011011001101" => rgb <= "111111";
            when "0011011001110" => rgb <= "111111";
            when "0011011001111" => rgb <= "111111";
            when "0011011010000" => rgb <= "000000";
            when "0011011010001" => rgb <= "000000";
            when "0011011010010" => rgb <= "111111";
            when "0011011010011" => rgb <= "111111";
            when "0011011010100" => rgb <= "111111";
            when "0011011010101" => rgb <= "111111";
            when "0011011010110" => rgb <= "111111";
            when "0011011010111" => rgb <= "111111";
            when "0011011011000" => rgb <= "000000";
            when "0011011011001" => rgb <= "000000";
            when "0011011011010" => rgb <= "111111";
            when "0011011011011" => rgb <= "111111";
            when "0011011011100" => rgb <= "111111";
            when "0011011011101" => rgb <= "111111";
            when "0011011011110" => rgb <= "111111";
            when "0011011011111" => rgb <= "111111";
            when "0011011100000" => rgb <= "111111";
            when "0011011100001" => rgb <= "010101";
            when "0011011100010" => rgb <= "100001";
            when "0011011100011" => rgb <= "100001";
            when "0011011100100" => rgb <= "100001";
            when "0011011100101" => rgb <= "100001";
            when "0011011100110" => rgb <= "100001";
            when "0011011100111" => rgb <= "100001";
            when "0011100000000" => rgb <= "100001";
            when "0011100000001" => rgb <= "100001";
            when "0011100000010" => rgb <= "100001";
            when "0011100000011" => rgb <= "100001";
            when "0011100000100" => rgb <= "100001";
            when "0011100000101" => rgb <= "100001";
            when "0011100000110" => rgb <= "100001";
            when "0011100000111" => rgb <= "010101";
            when "0011100001000" => rgb <= "101010";
            when "0011100001001" => rgb <= "101010";
            when "0011100001010" => rgb <= "111111";
            when "0011100001011" => rgb <= "111111";
            when "0011100001100" => rgb <= "111111";
            when "0011100001101" => rgb <= "111111";
            when "0011100001110" => rgb <= "111111";
            when "0011100001111" => rgb <= "111111";
            when "0011100010000" => rgb <= "000000";
            when "0011100010001" => rgb <= "000000";
            when "0011100010010" => rgb <= "111111";
            when "0011100010011" => rgb <= "111111";
            when "0011100010100" => rgb <= "111111";
            when "0011100010101" => rgb <= "111111";
            when "0011100010110" => rgb <= "111111";
            when "0011100010111" => rgb <= "111111";
            when "0011100011000" => rgb <= "000000";
            when "0011100011001" => rgb <= "000000";
            when "0011100011010" => rgb <= "111111";
            when "0011100011011" => rgb <= "111111";
            when "0011100011100" => rgb <= "111111";
            when "0011100011101" => rgb <= "111111";
            when "0011100011110" => rgb <= "111111";
            when "0011100011111" => rgb <= "111111";
            when "0011100100000" => rgb <= "111111";
            when "0011100100001" => rgb <= "010101";
            when "0011100100010" => rgb <= "100001";
            when "0011100100011" => rgb <= "100001";
            when "0011100100100" => rgb <= "100001";
            when "0011100100101" => rgb <= "100001";
            when "0011100100110" => rgb <= "100001";
            when "0011100100111" => rgb <= "100001";
            when "0011101000000" => rgb <= "100001";
            when "0011101000001" => rgb <= "100001";
            when "0011101000010" => rgb <= "100001";
            when "0011101000011" => rgb <= "100001";
            when "0011101000100" => rgb <= "100001";
            when "0011101000101" => rgb <= "100001";
            when "0011101000110" => rgb <= "100001";
            when "0011101000111" => rgb <= "010101";
            when "0011101001000" => rgb <= "101010";
            when "0011101001001" => rgb <= "101010";
            when "0011101001010" => rgb <= "111111";
            when "0011101001011" => rgb <= "111111";
            when "0011101001100" => rgb <= "111111";
            when "0011101001101" => rgb <= "111111";
            when "0011101001110" => rgb <= "111111";
            when "0011101001111" => rgb <= "111111";
            when "0011101010000" => rgb <= "000000";
            when "0011101010001" => rgb <= "000000";
            when "0011101010010" => rgb <= "111111";
            when "0011101010011" => rgb <= "111111";
            when "0011101010100" => rgb <= "111111";
            when "0011101010101" => rgb <= "111111";
            when "0011101010110" => rgb <= "111111";
            when "0011101010111" => rgb <= "111111";
            when "0011101011000" => rgb <= "000000";
            when "0011101011001" => rgb <= "000000";
            when "0011101011010" => rgb <= "111111";
            when "0011101011011" => rgb <= "111111";
            when "0011101011100" => rgb <= "111111";
            when "0011101011101" => rgb <= "111111";
            when "0011101011110" => rgb <= "111111";
            when "0011101011111" => rgb <= "111111";
            when "0011101100000" => rgb <= "111111";
            when "0011101100001" => rgb <= "010101";
            when "0011101100010" => rgb <= "100001";
            when "0011101100011" => rgb <= "100001";
            when "0011101100100" => rgb <= "100001";
            when "0011101100101" => rgb <= "100001";
            when "0011101100110" => rgb <= "100001";
            when "0011101100111" => rgb <= "100001";
            when "0011110000000" => rgb <= "100001";
            when "0011110000001" => rgb <= "100001";
            when "0011110000010" => rgb <= "100001";
            when "0011110000011" => rgb <= "100001";
            when "0011110000100" => rgb <= "100001";
            when "0011110000101" => rgb <= "100001";
            when "0011110000110" => rgb <= "100001";
            when "0011110000111" => rgb <= "010101";
            when "0011110001000" => rgb <= "101010";
            when "0011110001001" => rgb <= "101010";
            when "0011110001010" => rgb <= "111111";
            when "0011110001011" => rgb <= "111111";
            when "0011110001100" => rgb <= "111111";
            when "0011110001101" => rgb <= "111111";
            when "0011110001110" => rgb <= "111111";
            when "0011110001111" => rgb <= "111111";
            when "0011110010000" => rgb <= "000000";
            when "0011110010001" => rgb <= "000000";
            when "0011110010010" => rgb <= "111111";
            when "0011110010011" => rgb <= "111111";
            when "0011110010100" => rgb <= "111111";
            when "0011110010101" => rgb <= "111111";
            when "0011110010110" => rgb <= "111111";
            when "0011110010111" => rgb <= "111111";
            when "0011110011000" => rgb <= "000000";
            when "0011110011001" => rgb <= "000000";
            when "0011110011010" => rgb <= "111111";
            when "0011110011011" => rgb <= "111111";
            when "0011110011100" => rgb <= "111111";
            when "0011110011101" => rgb <= "111111";
            when "0011110011110" => rgb <= "111111";
            when "0011110011111" => rgb <= "111111";
            when "0011110100000" => rgb <= "111111";
            when "0011110100001" => rgb <= "010101";
            when "0011110100010" => rgb <= "100001";
            when "0011110100011" => rgb <= "100001";
            when "0011110100100" => rgb <= "100001";
            when "0011110100101" => rgb <= "100001";
            when "0011110100110" => rgb <= "100001";
            when "0011110100111" => rgb <= "100001";
            when "0011111000000" => rgb <= "100001";
            when "0011111000001" => rgb <= "100001";
            when "0011111000010" => rgb <= "100001";
            when "0011111000011" => rgb <= "100001";
            when "0011111000100" => rgb <= "100001";
            when "0011111000101" => rgb <= "100001";
            when "0011111000110" => rgb <= "100001";
            when "0011111000111" => rgb <= "010101";
            when "0011111001000" => rgb <= "101010";
            when "0011111001001" => rgb <= "101010";
            when "0011111001010" => rgb <= "111111";
            when "0011111001011" => rgb <= "111111";
            when "0011111001100" => rgb <= "111111";
            when "0011111001101" => rgb <= "111111";
            when "0011111001110" => rgb <= "111111";
            when "0011111001111" => rgb <= "111111";
            when "0011111010000" => rgb <= "000000";
            when "0011111010001" => rgb <= "000000";
            when "0011111010010" => rgb <= "111111";
            when "0011111010011" => rgb <= "111111";
            when "0011111010100" => rgb <= "111111";
            when "0011111010101" => rgb <= "111111";
            when "0011111010110" => rgb <= "111111";
            when "0011111010111" => rgb <= "111111";
            when "0011111011000" => rgb <= "000000";
            when "0011111011001" => rgb <= "000000";
            when "0011111011010" => rgb <= "111111";
            when "0011111011011" => rgb <= "111111";
            when "0011111011100" => rgb <= "111111";
            when "0011111011101" => rgb <= "111111";
            when "0011111011110" => rgb <= "111111";
            when "0011111011111" => rgb <= "111111";
            when "0011111100000" => rgb <= "111111";
            when "0011111100001" => rgb <= "010101";
            when "0011111100010" => rgb <= "100001";
            when "0011111100011" => rgb <= "100001";
            when "0011111100100" => rgb <= "100001";
            when "0011111100101" => rgb <= "100001";
            when "0011111100110" => rgb <= "100001";
            when "0011111100111" => rgb <= "100001";
            when "0100000000000" => rgb <= "100001";
            when "0100000000001" => rgb <= "100001";
            when "0100000000010" => rgb <= "100001";
            when "0100000000011" => rgb <= "100001";
            when "0100000000100" => rgb <= "100001";
            when "0100000000101" => rgb <= "100001";
            when "0100000000110" => rgb <= "100001";
            when "0100000000111" => rgb <= "010101";
            when "0100000001000" => rgb <= "101010";
            when "0100000001001" => rgb <= "101010";
            when "0100000001010" => rgb <= "111111";
            when "0100000001011" => rgb <= "111111";
            when "0100000001100" => rgb <= "111111";
            when "0100000001101" => rgb <= "111111";
            when "0100000001110" => rgb <= "111111";
            when "0100000001111" => rgb <= "111111";
            when "0100000010000" => rgb <= "111111";
            when "0100000010001" => rgb <= "111111";
            when "0100000010010" => rgb <= "111111";
            when "0100000010011" => rgb <= "111111";
            when "0100000010100" => rgb <= "111111";
            when "0100000010101" => rgb <= "001011";
            when "0100000010110" => rgb <= "001011";
            when "0100000010111" => rgb <= "001011";
            when "0100000011000" => rgb <= "001011";
            when "0100000011001" => rgb <= "001011";
            when "0100000011010" => rgb <= "001011";
            when "0100000011011" => rgb <= "001011";
            when "0100000011100" => rgb <= "001011";
            when "0100000011101" => rgb <= "001011";
            when "0100000011110" => rgb <= "001011";
            when "0100000011111" => rgb <= "111111";
            when "0100000100000" => rgb <= "111111";
            when "0100000100001" => rgb <= "010101";
            when "0100000100010" => rgb <= "100001";
            when "0100000100011" => rgb <= "100001";
            when "0100000100100" => rgb <= "100001";
            when "0100000100101" => rgb <= "100001";
            when "0100000100110" => rgb <= "100001";
            when "0100000100111" => rgb <= "100001";
            when "0100001000000" => rgb <= "100001";
            when "0100001000001" => rgb <= "100001";
            when "0100001000010" => rgb <= "100001";
            when "0100001000011" => rgb <= "100001";
            when "0100001000100" => rgb <= "100001";
            when "0100001000101" => rgb <= "100001";
            when "0100001000110" => rgb <= "100001";
            when "0100001000111" => rgb <= "010101";
            when "0100001001000" => rgb <= "101010";
            when "0100001001001" => rgb <= "101010";
            when "0100001001010" => rgb <= "111111";
            when "0100001001011" => rgb <= "111111";
            when "0100001001100" => rgb <= "111111";
            when "0100001001101" => rgb <= "111111";
            when "0100001001110" => rgb <= "111111";
            when "0100001001111" => rgb <= "111111";
            when "0100001010000" => rgb <= "111111";
            when "0100001010001" => rgb <= "111111";
            when "0100001010010" => rgb <= "111111";
            when "0100001010011" => rgb <= "111111";
            when "0100001010100" => rgb <= "111111";
            when "0100001010101" => rgb <= "001011";
            when "0100001010110" => rgb <= "001011";
            when "0100001010111" => rgb <= "001011";
            when "0100001011000" => rgb <= "001011";
            when "0100001011001" => rgb <= "001011";
            when "0100001011010" => rgb <= "001011";
            when "0100001011011" => rgb <= "001011";
            when "0100001011100" => rgb <= "001011";
            when "0100001011101" => rgb <= "001011";
            when "0100001011110" => rgb <= "001011";
            when "0100001011111" => rgb <= "111111";
            when "0100001100000" => rgb <= "111111";
            when "0100001100001" => rgb <= "010101";
            when "0100001100010" => rgb <= "100001";
            when "0100001100011" => rgb <= "100001";
            when "0100001100100" => rgb <= "100001";
            when "0100001100101" => rgb <= "100001";
            when "0100001100110" => rgb <= "100001";
            when "0100001100111" => rgb <= "100001";
            when "0100010000000" => rgb <= "100001";
            when "0100010000001" => rgb <= "100001";
            when "0100010000010" => rgb <= "100001";
            when "0100010000011" => rgb <= "100001";
            when "0100010000100" => rgb <= "100001";
            when "0100010000101" => rgb <= "100001";
            when "0100010000110" => rgb <= "100001";
            when "0100010000111" => rgb <= "010101";
            when "0100010001000" => rgb <= "101010";
            when "0100010001001" => rgb <= "101010";
            when "0100010001010" => rgb <= "111111";
            when "0100010001011" => rgb <= "111111";
            when "0100010001100" => rgb <= "111111";
            when "0100010001101" => rgb <= "111111";
            when "0100010001110" => rgb <= "111111";
            when "0100010001111" => rgb <= "111111";
            when "0100010010000" => rgb <= "111111";
            when "0100010010001" => rgb <= "111111";
            when "0100010010010" => rgb <= "111111";
            when "0100010010011" => rgb <= "111111";
            when "0100010010100" => rgb <= "111111";
            when "0100010010101" => rgb <= "001011";
            when "0100010010110" => rgb <= "001011";
            when "0100010010111" => rgb <= "001011";
            when "0100010011000" => rgb <= "001011";
            when "0100010011001" => rgb <= "001011";
            when "0100010011010" => rgb <= "001011";
            when "0100010011011" => rgb <= "001011";
            when "0100010011100" => rgb <= "001011";
            when "0100010011101" => rgb <= "001011";
            when "0100010011110" => rgb <= "001011";
            when "0100010011111" => rgb <= "111111";
            when "0100010100000" => rgb <= "111111";
            when "0100010100001" => rgb <= "010101";
            when "0100010100010" => rgb <= "100001";
            when "0100010100011" => rgb <= "100001";
            when "0100010100100" => rgb <= "100001";
            when "0100010100101" => rgb <= "100001";
            when "0100010100110" => rgb <= "100001";
            when "0100010100111" => rgb <= "100001";
            when "0100011000000" => rgb <= "100001";
            when "0100011000001" => rgb <= "100001";
            when "0100011000010" => rgb <= "000110";
            when "0100011000011" => rgb <= "100001";
            when "0100011000100" => rgb <= "100001";
            when "0100011000101" => rgb <= "100001";
            when "0100011000110" => rgb <= "100001";
            when "0100011000111" => rgb <= "100001";
            when "0100011001000" => rgb <= "010101";
            when "0100011001001" => rgb <= "101010";
            when "0100011001010" => rgb <= "111111";
            when "0100011001011" => rgb <= "111111";
            when "0100011001100" => rgb <= "111111";
            when "0100011001101" => rgb <= "111111";
            when "0100011001110" => rgb <= "111111";
            when "0100011001111" => rgb <= "111111";
            when "0100011010000" => rgb <= "111111";
            when "0100011010001" => rgb <= "111111";
            when "0100011010010" => rgb <= "111111";
            when "0100011010011" => rgb <= "111111";
            when "0100011010100" => rgb <= "111111";
            when "0100011010101" => rgb <= "111111";
            when "0100011010110" => rgb <= "111111";
            when "0100011010111" => rgb <= "111111";
            when "0100011011000" => rgb <= "111111";
            when "0100011011001" => rgb <= "111111";
            when "0100011011010" => rgb <= "111111";
            when "0100011011011" => rgb <= "111111";
            when "0100011011100" => rgb <= "111111";
            when "0100011011101" => rgb <= "111111";
            when "0100011011110" => rgb <= "111111";
            when "0100011011111" => rgb <= "111111";
            when "0100011100000" => rgb <= "010101";
            when "0100011100001" => rgb <= "100001";
            when "0100011100010" => rgb <= "100001";
            when "0100011100011" => rgb <= "100001";
            when "0100011100100" => rgb <= "100001";
            when "0100011100101" => rgb <= "100001";
            when "0100011100110" => rgb <= "100001";
            when "0100011100111" => rgb <= "100001";
            when "0100100000000" => rgb <= "100001";
            when "0100100000001" => rgb <= "100001";
            when "0100100000010" => rgb <= "100001";
            when "0100100000011" => rgb <= "000110";
            when "0100100000100" => rgb <= "100001";
            when "0100100000101" => rgb <= "100001";
            when "0100100000110" => rgb <= "000110";
            when "0100100000111" => rgb <= "100001";
            when "0100100001000" => rgb <= "010101";
            when "0100100001001" => rgb <= "101010";
            when "0100100001010" => rgb <= "101010";
            when "0100100001011" => rgb <= "111111";
            when "0100100001100" => rgb <= "111111";
            when "0100100001101" => rgb <= "111111";
            when "0100100001110" => rgb <= "111111";
            when "0100100001111" => rgb <= "111111";
            when "0100100010000" => rgb <= "111111";
            when "0100100010001" => rgb <= "111111";
            when "0100100010010" => rgb <= "111111";
            when "0100100010011" => rgb <= "111111";
            when "0100100010100" => rgb <= "111111";
            when "0100100010101" => rgb <= "111111";
            when "0100100010110" => rgb <= "111111";
            when "0100100010111" => rgb <= "111111";
            when "0100100011000" => rgb <= "111111";
            when "0100100011001" => rgb <= "111111";
            when "0100100011010" => rgb <= "111111";
            when "0100100011011" => rgb <= "111111";
            when "0100100011100" => rgb <= "111111";
            when "0100100011101" => rgb <= "111111";
            when "0100100011110" => rgb <= "111111";
            when "0100100011111" => rgb <= "111111";
            when "0100100100000" => rgb <= "010101";
            when "0100100100001" => rgb <= "100001";
            when "0100100100010" => rgb <= "100001";
            when "0100100100011" => rgb <= "100001";
            when "0100100100100" => rgb <= "100001";
            when "0100100100101" => rgb <= "100001";
            when "0100100100110" => rgb <= "100001";
            when "0100100100111" => rgb <= "100001";
            when "0100101000000" => rgb <= "100001";
            when "0100101000001" => rgb <= "100001";
            when "0100101000010" => rgb <= "100001";
            when "0100101000011" => rgb <= "000110";
            when "0100101000100" => rgb <= "100001";
            when "0100101000101" => rgb <= "000110";
            when "0100101000110" => rgb <= "100001";
            when "0100101000111" => rgb <= "100001";
            when "0100101001000" => rgb <= "100001";
            when "0100101001001" => rgb <= "010101";
            when "0100101001010" => rgb <= "101010";
            when "0100101001011" => rgb <= "101010";
            when "0100101001100" => rgb <= "111111";
            when "0100101001101" => rgb <= "111111";
            when "0100101001110" => rgb <= "111111";
            when "0100101001111" => rgb <= "111111";
            when "0100101010000" => rgb <= "111111";
            when "0100101010001" => rgb <= "111111";
            when "0100101010010" => rgb <= "111111";
            when "0100101010011" => rgb <= "111111";
            when "0100101010100" => rgb <= "111111";
            when "0100101010101" => rgb <= "111111";
            when "0100101010110" => rgb <= "111111";
            when "0100101010111" => rgb <= "111111";
            when "0100101011000" => rgb <= "111111";
            when "0100101011001" => rgb <= "111111";
            when "0100101011010" => rgb <= "111111";
            when "0100101011011" => rgb <= "111111";
            when "0100101011100" => rgb <= "111111";
            when "0100101011101" => rgb <= "111111";
            when "0100101011110" => rgb <= "111111";
            when "0100101011111" => rgb <= "010101";
            when "0100101100000" => rgb <= "100001";
            when "0100101100001" => rgb <= "100001";
            when "0100101100010" => rgb <= "000110";
            when "0100101100011" => rgb <= "100001";
            when "0100101100100" => rgb <= "100001";
            when "0100101100101" => rgb <= "000110";
            when "0100101100110" => rgb <= "100001";
            when "0100101100111" => rgb <= "100001";
            when "0100110000000" => rgb <= "100001";
            when "0100110000001" => rgb <= "100001";
            when "0100110000010" => rgb <= "100001";
            when "0100110000011" => rgb <= "000110";
            when "0100110000100" => rgb <= "100001";
            when "0100110000101" => rgb <= "000110";
            when "0100110000110" => rgb <= "100001";
            when "0100110000111" => rgb <= "100001";
            when "0100110001000" => rgb <= "100001";
            when "0100110001001" => rgb <= "010101";
            when "0100110001010" => rgb <= "101010";
            when "0100110001011" => rgb <= "101010";
            when "0100110001100" => rgb <= "111111";
            when "0100110001101" => rgb <= "111111";
            when "0100110001110" => rgb <= "111111";
            when "0100110001111" => rgb <= "111111";
            when "0100110010000" => rgb <= "111111";
            when "0100110010001" => rgb <= "111111";
            when "0100110010010" => rgb <= "111111";
            when "0100110010011" => rgb <= "111111";
            when "0100110010100" => rgb <= "111111";
            when "0100110010101" => rgb <= "111111";
            when "0100110010110" => rgb <= "111111";
            when "0100110010111" => rgb <= "111111";
            when "0100110011000" => rgb <= "111111";
            when "0100110011001" => rgb <= "111111";
            when "0100110011010" => rgb <= "111111";
            when "0100110011011" => rgb <= "111111";
            when "0100110011100" => rgb <= "111111";
            when "0100110011101" => rgb <= "111111";
            when "0100110011110" => rgb <= "111111";
            when "0100110011111" => rgb <= "010101";
            when "0100110100000" => rgb <= "100001";
            when "0100110100001" => rgb <= "100001";
            when "0100110100010" => rgb <= "000110";
            when "0100110100011" => rgb <= "100001";
            when "0100110100100" => rgb <= "100001";
            when "0100110100101" => rgb <= "000110";
            when "0100110100110" => rgb <= "100001";
            when "0100110100111" => rgb <= "100001";
            when "0100111000000" => rgb <= "000110";
            when "0100111000001" => rgb <= "000110";
            when "0100111000010" => rgb <= "100001";
            when "0100111000011" => rgb <= "100001";
            when "0100111000100" => rgb <= "000110";
            when "0100111000101" => rgb <= "000110";
            when "0100111000110" => rgb <= "100001";
            when "0100111000111" => rgb <= "100001";
            when "0100111001000" => rgb <= "100001";
            when "0100111001001" => rgb <= "100001";
            when "0100111001010" => rgb <= "010101";
            when "0100111001011" => rgb <= "101010";
            when "0100111001100" => rgb <= "101010";
            when "0100111001101" => rgb <= "111111";
            when "0100111001110" => rgb <= "111111";
            when "0100111001111" => rgb <= "111111";
            when "0100111010000" => rgb <= "111111";
            when "0100111010001" => rgb <= "111111";
            when "0100111010010" => rgb <= "111111";
            when "0100111010011" => rgb <= "111111";
            when "0100111010100" => rgb <= "111111";
            when "0100111010101" => rgb <= "111111";
            when "0100111010110" => rgb <= "111111";
            when "0100111010111" => rgb <= "111111";
            when "0100111011000" => rgb <= "111111";
            when "0100111011001" => rgb <= "111111";
            when "0100111011010" => rgb <= "111111";
            when "0100111011011" => rgb <= "111111";
            when "0100111011100" => rgb <= "111111";
            when "0100111011101" => rgb <= "111111";
            when "0100111011110" => rgb <= "010101";
            when "0100111011111" => rgb <= "100001";
            when "0100111100000" => rgb <= "100001";
            when "0100111100001" => rgb <= "100001";
            when "0100111100010" => rgb <= "000110";
            when "0100111100011" => rgb <= "100001";
            when "0100111100100" => rgb <= "000110";
            when "0100111100101" => rgb <= "100001";
            when "0100111100110" => rgb <= "100001";
            when "0100111100111" => rgb <= "100001";
            when "0101000000000" => rgb <= "100001";
            when "0101000000001" => rgb <= "100001";
            when "0101000000010" => rgb <= "000110";
            when "0101000000011" => rgb <= "000110";
            when "0101000000100" => rgb <= "000110";
            when "0101000000101" => rgb <= "100001";
            when "0101000000110" => rgb <= "100001";
            when "0101000000111" => rgb <= "000001";
            when "0101000001000" => rgb <= "000001";
            when "0101000001001" => rgb <= "000010";
            when "0101000001010" => rgb <= "000010";
            when "0101000001011" => rgb <= "000010";
            when "0101000001100" => rgb <= "000010";
            when "0101000001101" => rgb <= "000010";
            when "0101000001110" => rgb <= "000010";
            when "0101000001111" => rgb <= "000010";
            when "0101000010000" => rgb <= "000010";
            when "0101000010001" => rgb <= "000010";
            when "0101000010010" => rgb <= "000010";
            when "0101000010011" => rgb <= "000010";
            when "0101000010100" => rgb <= "000010";
            when "0101000010101" => rgb <= "000010";
            when "0101000010110" => rgb <= "000010";
            when "0101000010111" => rgb <= "000010";
            when "0101000011000" => rgb <= "000010";
            when "0101000011001" => rgb <= "000010";
            when "0101000011010" => rgb <= "000010";
            when "0101000011011" => rgb <= "000010";
            when "0101000011100" => rgb <= "000010";
            when "0101000011101" => rgb <= "000001";
            when "0101000011110" => rgb <= "000001";
            when "0101000011111" => rgb <= "100001";
            when "0101000100000" => rgb <= "100001";
            when "0101000100001" => rgb <= "100001";
            when "0101000100010" => rgb <= "100001";
            when "0101000100011" => rgb <= "000110";
            when "0101000100100" => rgb <= "100001";
            when "0101000100101" => rgb <= "100001";
            when "0101000100110" => rgb <= "100001";
            when "0101000100111" => rgb <= "100001";
            when "0101001000000" => rgb <= "100001";
            when "0101001000001" => rgb <= "100001";
            when "0101001000010" => rgb <= "100001";
            when "0101001000011" => rgb <= "100001";
            when "0101001000100" => rgb <= "000110";
            when "0101001000101" => rgb <= "000110";
            when "0101001000110" => rgb <= "100001";
            when "0101001000111" => rgb <= "000001";
            when "0101001001000" => rgb <= "000010";
            when "0101001001001" => rgb <= "000010";
            when "0101001001010" => rgb <= "000010";
            when "0101001001011" => rgb <= "000010";
            when "0101001001100" => rgb <= "000010";
            when "0101001001101" => rgb <= "000010";
            when "0101001001110" => rgb <= "000010";
            when "0101001001111" => rgb <= "000010";
            when "0101001010000" => rgb <= "000010";
            when "0101001010001" => rgb <= "000010";
            when "0101001010010" => rgb <= "000010";
            when "0101001010011" => rgb <= "000010";
            when "0101001010100" => rgb <= "000010";
            when "0101001010101" => rgb <= "000010";
            when "0101001010110" => rgb <= "000010";
            when "0101001010111" => rgb <= "000010";
            when "0101001011000" => rgb <= "000010";
            when "0101001011001" => rgb <= "000010";
            when "0101001011010" => rgb <= "000010";
            when "0101001011011" => rgb <= "000010";
            when "0101001011100" => rgb <= "000010";
            when "0101001011101" => rgb <= "000001";
            when "0101001011110" => rgb <= "000001";
            when "0101001011111" => rgb <= "100001";
            when "0101001100000" => rgb <= "100001";
            when "0101001100001" => rgb <= "100001";
            when "0101001100010" => rgb <= "100001";
            when "0101001100011" => rgb <= "000110";
            when "0101001100100" => rgb <= "000110";
            when "0101001100101" => rgb <= "100001";
            when "0101001100110" => rgb <= "000110";
            when "0101001100111" => rgb <= "000110";
            when "0101010000000" => rgb <= "100001";
            when "0101010000001" => rgb <= "100001";
            when "0101010000010" => rgb <= "100001";
            when "0101010000011" => rgb <= "100001";
            when "0101010000100" => rgb <= "000110";
            when "0101010000101" => rgb <= "000110";
            when "0101010000110" => rgb <= "100001";
            when "0101010000111" => rgb <= "000001";
            when "0101010001000" => rgb <= "000010";
            when "0101010001001" => rgb <= "000010";
            when "0101010001010" => rgb <= "000010";
            when "0101010001011" => rgb <= "000010";
            when "0101010001100" => rgb <= "000010";
            when "0101010001101" => rgb <= "000010";
            when "0101010001110" => rgb <= "000010";
            when "0101010001111" => rgb <= "000010";
            when "0101010010000" => rgb <= "000010";
            when "0101010010001" => rgb <= "000010";
            when "0101010010010" => rgb <= "000010";
            when "0101010010011" => rgb <= "000010";
            when "0101010010100" => rgb <= "000010";
            when "0101010010101" => rgb <= "000010";
            when "0101010010110" => rgb <= "000010";
            when "0101010010111" => rgb <= "000010";
            when "0101010011000" => rgb <= "000010";
            when "0101010011001" => rgb <= "000010";
            when "0101010011010" => rgb <= "000010";
            when "0101010011011" => rgb <= "000010";
            when "0101010011100" => rgb <= "000010";
            when "0101010011101" => rgb <= "000001";
            when "0101010011110" => rgb <= "000001";
            when "0101010011111" => rgb <= "100001";
            when "0101010100000" => rgb <= "100001";
            when "0101010100001" => rgb <= "100001";
            when "0101010100010" => rgb <= "100001";
            when "0101010100011" => rgb <= "000110";
            when "0101010100100" => rgb <= "000110";
            when "0101010100101" => rgb <= "100001";
            when "0101010100110" => rgb <= "000110";
            when "0101010100111" => rgb <= "000110";
            when "0101011000000" => rgb <= "100001";
            when "0101011000001" => rgb <= "100001";
            when "0101011000010" => rgb <= "100001";
            when "0101011000011" => rgb <= "100001";
            when "0101011000100" => rgb <= "100001";
            when "0101011000101" => rgb <= "000110";
            when "0101011000110" => rgb <= "000110";
            when "0101011000111" => rgb <= "000010";
            when "0101011001000" => rgb <= "000010";
            when "0101011001001" => rgb <= "000010";
            when "0101011001010" => rgb <= "000010";
            when "0101011001011" => rgb <= "000010";
            when "0101011001100" => rgb <= "000010";
            when "0101011001101" => rgb <= "000010";
            when "0101011001110" => rgb <= "000010";
            when "0101011001111" => rgb <= "000010";
            when "0101011010000" => rgb <= "000010";
            when "0101011010001" => rgb <= "000010";
            when "0101011010010" => rgb <= "000010";
            when "0101011010011" => rgb <= "000010";
            when "0101011010100" => rgb <= "000010";
            when "0101011010101" => rgb <= "000010";
            when "0101011010110" => rgb <= "000010";
            when "0101011010111" => rgb <= "000010";
            when "0101011011000" => rgb <= "000010";
            when "0101011011001" => rgb <= "000010";
            when "0101011011010" => rgb <= "000010";
            when "0101011011011" => rgb <= "000010";
            when "0101011011100" => rgb <= "000010";
            when "0101011011101" => rgb <= "000001";
            when "0101011011110" => rgb <= "000001";
            when "0101011011111" => rgb <= "010101";
            when "0101011100000" => rgb <= "100001";
            when "0101011100001" => rgb <= "100001";
            when "0101011100010" => rgb <= "100001";
            when "0101011100011" => rgb <= "000110";
            when "0101011100100" => rgb <= "000110";
            when "0101011100101" => rgb <= "000110";
            when "0101011100110" => rgb <= "100001";
            when "0101011100111" => rgb <= "100001";
            when "0101100000000" => rgb <= "100001";
            when "0101100000001" => rgb <= "100001";
            when "0101100000010" => rgb <= "100001";
            when "0101100000011" => rgb <= "100001";
            when "0101100000100" => rgb <= "100001";
            when "0101100000101" => rgb <= "000001";
            when "0101100000110" => rgb <= "000110";
            when "0101100000111" => rgb <= "000110";
            when "0101100001000" => rgb <= "000010";
            when "0101100001001" => rgb <= "010101";
            when "0101100001010" => rgb <= "010101";
            when "0101100001011" => rgb <= "010101";
            when "0101100001100" => rgb <= "101010";
            when "0101100001101" => rgb <= "101010";
            when "0101100001110" => rgb <= "111111";
            when "0101100001111" => rgb <= "111111";
            when "0101100010000" => rgb <= "111111";
            when "0101100010001" => rgb <= "111111";
            when "0101100010010" => rgb <= "111111";
            when "0101100010011" => rgb <= "111111";
            when "0101100010100" => rgb <= "111111";
            when "0101100010101" => rgb <= "111111";
            when "0101100010110" => rgb <= "111111";
            when "0101100010111" => rgb <= "111111";
            when "0101100011000" => rgb <= "111111";
            when "0101100011001" => rgb <= "111111";
            when "0101100011010" => rgb <= "111111";
            when "0101100011011" => rgb <= "111111";
            when "0101100011100" => rgb <= "111111";
            when "0101100011101" => rgb <= "111111";
            when "0101100011110" => rgb <= "111111";
            when "0101100011111" => rgb <= "111111";
            when "0101100100000" => rgb <= "010101";
            when "0101100100001" => rgb <= "100001";
            when "0101100100010" => rgb <= "000110";
            when "0101100100011" => rgb <= "000110";
            when "0101100100100" => rgb <= "100001";
            when "0101100100101" => rgb <= "100001";
            when "0101100100110" => rgb <= "100001";
            when "0101100100111" => rgb <= "100001";
            when "0101101000000" => rgb <= "100001";
            when "0101101000001" => rgb <= "100001";
            when "0101101000010" => rgb <= "100001";
            when "0101101000011" => rgb <= "100001";
            when "0101101000100" => rgb <= "000001";
            when "0101101000101" => rgb <= "000001";
            when "0101101000110" => rgb <= "000010";
            when "0101101000111" => rgb <= "000110";
            when "0101101001000" => rgb <= "000110";
            when "0101101001001" => rgb <= "010101";
            when "0101101001010" => rgb <= "101010";
            when "0101101001011" => rgb <= "101010";
            when "0101101001100" => rgb <= "101010";
            when "0101101001101" => rgb <= "111111";
            when "0101101001110" => rgb <= "111111";
            when "0101101001111" => rgb <= "111111";
            when "0101101010000" => rgb <= "111111";
            when "0101101010001" => rgb <= "111111";
            when "0101101010010" => rgb <= "111111";
            when "0101101010011" => rgb <= "111111";
            when "0101101010100" => rgb <= "111111";
            when "0101101010101" => rgb <= "111111";
            when "0101101010110" => rgb <= "111111";
            when "0101101010111" => rgb <= "111111";
            when "0101101011000" => rgb <= "111111";
            when "0101101011001" => rgb <= "111111";
            when "0101101011010" => rgb <= "111111";
            when "0101101011011" => rgb <= "111111";
            when "0101101011100" => rgb <= "111111";
            when "0101101011101" => rgb <= "111111";
            when "0101101011110" => rgb <= "111111";
            when "0101101011111" => rgb <= "111111";
            when "0101101100000" => rgb <= "111111";
            when "0101101100001" => rgb <= "000110";
            when "0101101100010" => rgb <= "000110";
            when "0101101100011" => rgb <= "100001";
            when "0101101100100" => rgb <= "100001";
            when "0101101100101" => rgb <= "100001";
            when "0101101100110" => rgb <= "100001";
            when "0101101100111" => rgb <= "100001";
            when "0101110000000" => rgb <= "100001";
            when "0101110000001" => rgb <= "100001";
            when "0101110000010" => rgb <= "100001";
            when "0101110000011" => rgb <= "100001";
            when "0101110000100" => rgb <= "000001";
            when "0101110000101" => rgb <= "000001";
            when "0101110000110" => rgb <= "000010";
            when "0101110000111" => rgb <= "000110";
            when "0101110001000" => rgb <= "000110";
            when "0101110001001" => rgb <= "010101";
            when "0101110001010" => rgb <= "101010";
            when "0101110001011" => rgb <= "101010";
            when "0101110001100" => rgb <= "101010";
            when "0101110001101" => rgb <= "111111";
            when "0101110001110" => rgb <= "111111";
            when "0101110001111" => rgb <= "111111";
            when "0101110010000" => rgb <= "111111";
            when "0101110010001" => rgb <= "111111";
            when "0101110010010" => rgb <= "111111";
            when "0101110010011" => rgb <= "111111";
            when "0101110010100" => rgb <= "111111";
            when "0101110010101" => rgb <= "111111";
            when "0101110010110" => rgb <= "111111";
            when "0101110010111" => rgb <= "111111";
            when "0101110011000" => rgb <= "111111";
            when "0101110011001" => rgb <= "111111";
            when "0101110011010" => rgb <= "111111";
            when "0101110011011" => rgb <= "111111";
            when "0101110011100" => rgb <= "111111";
            when "0101110011101" => rgb <= "111111";
            when "0101110011110" => rgb <= "111111";
            when "0101110011111" => rgb <= "111111";
            when "0101110100000" => rgb <= "111111";
            when "0101110100001" => rgb <= "000110";
            when "0101110100010" => rgb <= "000110";
            when "0101110100011" => rgb <= "100001";
            when "0101110100100" => rgb <= "100001";
            when "0101110100101" => rgb <= "100001";
            when "0101110100110" => rgb <= "100001";
            when "0101110100111" => rgb <= "100001";
            when "0101111000000" => rgb <= "100001";
            when "0101111000001" => rgb <= "100001";
            when "0101111000010" => rgb <= "100001";
            when "0101111000011" => rgb <= "000001";
            when "0101111000100" => rgb <= "000001";
            when "0101111000101" => rgb <= "000010";
            when "0101111000110" => rgb <= "000010";
            when "0101111000111" => rgb <= "100001";
            when "0101111001000" => rgb <= "000110";
            when "0101111001001" => rgb <= "000110";
            when "0101111001010" => rgb <= "101010";
            when "0101111001011" => rgb <= "101010";
            when "0101111001100" => rgb <= "111111";
            when "0101111001101" => rgb <= "111111";
            when "0101111001110" => rgb <= "111111";
            when "0101111001111" => rgb <= "111111";
            when "0101111010000" => rgb <= "111111";
            when "0101111010001" => rgb <= "111111";
            when "0101111010010" => rgb <= "111111";
            when "0101111010011" => rgb <= "111111";
            when "0101111010100" => rgb <= "111111";
            when "0101111010101" => rgb <= "111111";
            when "0101111010110" => rgb <= "111111";
            when "0101111010111" => rgb <= "111111";
            when "0101111011000" => rgb <= "111111";
            when "0101111011001" => rgb <= "111111";
            when "0101111011010" => rgb <= "111111";
            when "0101111011011" => rgb <= "111111";
            when "0101111011100" => rgb <= "111111";
            when "0101111011101" => rgb <= "111111";
            when "0101111011110" => rgb <= "111111";
            when "0101111011111" => rgb <= "111111";
            when "0101111100000" => rgb <= "000110";
            when "0101111100001" => rgb <= "000110";
            when "0101111100010" => rgb <= "100001";
            when "0101111100011" => rgb <= "100001";
            when "0101111100100" => rgb <= "100001";
            when "0101111100101" => rgb <= "100001";
            when "0101111100110" => rgb <= "100001";
            when "0101111100111" => rgb <= "100001";
            when "0110000000000" => rgb <= "100001";
            when "0110000000001" => rgb <= "100001";
            when "0110000000010" => rgb <= "100001";
            when "0110000000011" => rgb <= "100001";
            when "0110000000100" => rgb <= "000010";
            when "0110000000101" => rgb <= "000010";
            when "0110000000110" => rgb <= "000010";
            when "0110000000111" => rgb <= "100001";
            when "0110000001000" => rgb <= "010101";
            when "0110000001001" => rgb <= "000110";
            when "0110000001010" => rgb <= "000110";
            when "0110000001011" => rgb <= "101010";
            when "0110000001100" => rgb <= "111111";
            when "0110000001101" => rgb <= "111111";
            when "0110000001110" => rgb <= "111111";
            when "0110000001111" => rgb <= "111111";
            when "0110000010000" => rgb <= "111111";
            when "0110000010001" => rgb <= "111111";
            when "0110000010010" => rgb <= "111111";
            when "0110000010011" => rgb <= "111111";
            when "0110000010100" => rgb <= "111111";
            when "0110000010101" => rgb <= "111111";
            when "0110000010110" => rgb <= "111111";
            when "0110000010111" => rgb <= "111111";
            when "0110000011000" => rgb <= "111111";
            when "0110000011001" => rgb <= "111111";
            when "0110000011010" => rgb <= "111111";
            when "0110000011011" => rgb <= "111111";
            when "0110000011100" => rgb <= "111111";
            when "0110000011101" => rgb <= "111111";
            when "0110000011110" => rgb <= "111111";
            when "0110000011111" => rgb <= "000110";
            when "0110000100000" => rgb <= "000110";
            when "0110000100001" => rgb <= "010101";
            when "0110000100010" => rgb <= "100001";
            when "0110000100011" => rgb <= "100001";
            when "0110000100100" => rgb <= "100001";
            when "0110000100101" => rgb <= "100001";
            when "0110000100110" => rgb <= "100001";
            when "0110000100111" => rgb <= "100001";
            when "0110001000000" => rgb <= "100001";
            when "0110001000001" => rgb <= "100001";
            when "0110001000010" => rgb <= "100001";
            when "0110001000011" => rgb <= "100001";
            when "0110001000100" => rgb <= "000010";
            when "0110001000101" => rgb <= "000010";
            when "0110001000110" => rgb <= "000010";
            when "0110001000111" => rgb <= "010101";
            when "0110001001000" => rgb <= "010101";
            when "0110001001001" => rgb <= "101010";
            when "0110001001010" => rgb <= "000110";
            when "0110001001011" => rgb <= "000110";
            when "0110001001100" => rgb <= "111111";
            when "0110001001101" => rgb <= "111111";
            when "0110001001110" => rgb <= "111111";
            when "0110001001111" => rgb <= "111111";
            when "0110001010000" => rgb <= "111111";
            when "0110001010001" => rgb <= "111111";
            when "0110001010010" => rgb <= "111111";
            when "0110001010011" => rgb <= "111111";
            when "0110001010100" => rgb <= "111111";
            when "0110001010101" => rgb <= "111111";
            when "0110001010110" => rgb <= "111111";
            when "0110001010111" => rgb <= "111111";
            when "0110001011000" => rgb <= "111111";
            when "0110001011001" => rgb <= "111111";
            when "0110001011010" => rgb <= "111111";
            when "0110001011011" => rgb <= "111111";
            when "0110001011100" => rgb <= "111111";
            when "0110001011101" => rgb <= "111111";
            when "0110001011110" => rgb <= "111111";
            when "0110001011111" => rgb <= "111111";
            when "0110001100000" => rgb <= "111111";
            when "0110001100001" => rgb <= "010101";
            when "0110001100010" => rgb <= "100001";
            when "0110001100011" => rgb <= "100001";
            when "0110001100100" => rgb <= "100001";
            when "0110001100101" => rgb <= "100001";
            when "0110001100110" => rgb <= "100001";
            when "0110001100111" => rgb <= "100001";
            when "0110010000000" => rgb <= "100001";
            when "0110010000001" => rgb <= "100001";
            when "0110010000010" => rgb <= "100001";
            when "0110010000011" => rgb <= "100001";
            when "0110010000100" => rgb <= "000010";
            when "0110010000101" => rgb <= "000010";
            when "0110010000110" => rgb <= "100001";
            when "0110010000111" => rgb <= "010101";
            when "0110010001000" => rgb <= "010101";
            when "0110010001001" => rgb <= "101010";
            when "0110010001010" => rgb <= "101010";
            when "0110010001011" => rgb <= "111111";
            when "0110010001100" => rgb <= "111111";
            when "0110010001101" => rgb <= "111111";
            when "0110010001110" => rgb <= "111111";
            when "0110010001111" => rgb <= "111111";
            when "0110010010000" => rgb <= "111111";
            when "0110010010001" => rgb <= "111111";
            when "0110010010010" => rgb <= "111111";
            when "0110010010011" => rgb <= "111111";
            when "0110010010100" => rgb <= "111111";
            when "0110010010101" => rgb <= "111111";
            when "0110010010110" => rgb <= "111111";
            when "0110010010111" => rgb <= "111111";
            when "0110010011000" => rgb <= "111111";
            when "0110010011001" => rgb <= "111111";
            when "0110010011010" => rgb <= "111111";
            when "0110010011011" => rgb <= "111111";
            when "0110010011100" => rgb <= "111111";
            when "0110010011101" => rgb <= "111111";
            when "0110010011110" => rgb <= "111111";
            when "0110010011111" => rgb <= "111111";
            when "0110010100000" => rgb <= "111111";
            when "0110010100001" => rgb <= "010101";
            when "0110010100010" => rgb <= "100001";
            when "0110010100011" => rgb <= "100001";
            when "0110010100100" => rgb <= "100001";
            when "0110010100101" => rgb <= "100001";
            when "0110010100110" => rgb <= "100001";
            when "0110010100111" => rgb <= "100001";
            when "0110011000000" => rgb <= "100001";
            when "0110011000001" => rgb <= "100001";
            when "0110011000010" => rgb <= "100001";
            when "0110011000011" => rgb <= "100001";
            when "0110011000100" => rgb <= "000010";
            when "0110011000101" => rgb <= "000010";
            when "0110011000110" => rgb <= "100001";
            when "0110011000111" => rgb <= "010101";
            when "0110011001000" => rgb <= "010101";
            when "0110011001001" => rgb <= "101010";
            when "0110011001010" => rgb <= "101010";
            when "0110011001011" => rgb <= "111111";
            when "0110011001100" => rgb <= "111111";
            when "0110011001101" => rgb <= "111111";
            when "0110011001110" => rgb <= "111111";
            when "0110011001111" => rgb <= "111111";
            when "0110011010000" => rgb <= "111111";
            when "0110011010001" => rgb <= "111111";
            when "0110011010010" => rgb <= "111111";
            when "0110011010011" => rgb <= "111111";
            when "0110011010100" => rgb <= "111111";
            when "0110011010101" => rgb <= "111111";
            when "0110011010110" => rgb <= "111111";
            when "0110011010111" => rgb <= "111111";
            when "0110011011000" => rgb <= "111111";
            when "0110011011001" => rgb <= "111111";
            when "0110011011010" => rgb <= "111111";
            when "0110011011011" => rgb <= "111111";
            when "0110011011100" => rgb <= "111111";
            when "0110011011101" => rgb <= "111111";
            when "0110011011110" => rgb <= "111111";
            when "0110011011111" => rgb <= "111111";
            when "0110011100000" => rgb <= "111111";
            when "0110011100001" => rgb <= "010101";
            when "0110011100010" => rgb <= "100001";
            when "0110011100011" => rgb <= "100001";
            when "0110011100100" => rgb <= "100001";
            when "0110011100101" => rgb <= "100001";
            when "0110011100110" => rgb <= "100001";
            when "0110011100111" => rgb <= "100001";
            when "0110100000000" => rgb <= "100001";
            when "0110100000001" => rgb <= "100001";
            when "0110100000010" => rgb <= "100001";
            when "0110100000011" => rgb <= "100001";
            when "0110100000100" => rgb <= "000010";
            when "0110100000101" => rgb <= "000010";
            when "0110100000110" => rgb <= "100001";
            when "0110100000111" => rgb <= "010101";
            when "0110100001000" => rgb <= "010101";
            when "0110100001001" => rgb <= "101010";
            when "0110100001010" => rgb <= "101010";
            when "0110100001011" => rgb <= "111111";
            when "0110100001100" => rgb <= "111111";
            when "0110100001101" => rgb <= "111111";
            when "0110100001110" => rgb <= "111111";
            when "0110100001111" => rgb <= "111111";
            when "0110100010000" => rgb <= "111111";
            when "0110100010001" => rgb <= "111111";
            when "0110100010010" => rgb <= "111111";
            when "0110100010011" => rgb <= "111111";
            when "0110100010100" => rgb <= "111111";
            when "0110100010101" => rgb <= "111111";
            when "0110100010110" => rgb <= "111111";
            when "0110100010111" => rgb <= "111111";
            when "0110100011000" => rgb <= "111111";
            when "0110100011001" => rgb <= "111111";
            when "0110100011010" => rgb <= "111111";
            when "0110100011011" => rgb <= "111111";
            when "0110100011100" => rgb <= "111111";
            when "0110100011101" => rgb <= "111111";
            when "0110100011110" => rgb <= "111111";
            when "0110100011111" => rgb <= "111111";
            when "0110100100000" => rgb <= "111111";
            when "0110100100001" => rgb <= "010101";
            when "0110100100010" => rgb <= "100001";
            when "0110100100011" => rgb <= "100001";
            when "0110100100100" => rgb <= "100001";
            when "0110100100101" => rgb <= "100001";
            when "0110100100110" => rgb <= "100001";
            when "0110100100111" => rgb <= "100001";
            when "0110101000000" => rgb <= "100001";
            when "0110101000001" => rgb <= "100001";
            when "0110101000010" => rgb <= "100001";
            when "0110101000011" => rgb <= "100001";
            when "0110101000100" => rgb <= "100001";
            when "0110101000101" => rgb <= "100001";
            when "0110101000110" => rgb <= "100001";
            when "0110101000111" => rgb <= "010101";
            when "0110101001000" => rgb <= "010101";
            when "0110101001001" => rgb <= "101010";
            when "0110101001010" => rgb <= "101010";
            when "0110101001011" => rgb <= "111111";
            when "0110101001100" => rgb <= "111111";
            when "0110101001101" => rgb <= "111111";
            when "0110101001110" => rgb <= "111111";
            when "0110101001111" => rgb <= "111111";
            when "0110101010000" => rgb <= "111111";
            when "0110101010001" => rgb <= "111111";
            when "0110101010010" => rgb <= "111111";
            when "0110101010011" => rgb <= "111111";
            when "0110101010100" => rgb <= "111111";
            when "0110101010101" => rgb <= "111111";
            when "0110101010110" => rgb <= "111111";
            when "0110101010111" => rgb <= "111111";
            when "0110101011000" => rgb <= "111111";
            when "0110101011001" => rgb <= "111111";
            when "0110101011010" => rgb <= "111111";
            when "0110101011011" => rgb <= "111111";
            when "0110101011100" => rgb <= "111111";
            when "0110101011101" => rgb <= "111111";
            when "0110101011110" => rgb <= "111111";
            when "0110101011111" => rgb <= "111111";
            when "0110101100000" => rgb <= "111111";
            when "0110101100001" => rgb <= "010101";
            when "0110101100010" => rgb <= "100001";
            when "0110101100011" => rgb <= "100001";
            when "0110101100100" => rgb <= "100001";
            when "0110101100101" => rgb <= "100001";
            when "0110101100110" => rgb <= "100001";
            when "0110101100111" => rgb <= "100001";
            when "0110110000000" => rgb <= "100001";
            when "0110110000001" => rgb <= "100001";
            when "0110110000010" => rgb <= "100001";
            when "0110110000011" => rgb <= "100001";
            when "0110110000100" => rgb <= "100001";
            when "0110110000101" => rgb <= "100001";
            when "0110110000110" => rgb <= "100001";
            when "0110110000111" => rgb <= "010101";
            when "0110110001000" => rgb <= "101010";
            when "0110110001001" => rgb <= "101010";
            when "0110110001010" => rgb <= "101010";
            when "0110110001011" => rgb <= "111111";
            when "0110110001100" => rgb <= "111111";
            when "0110110001101" => rgb <= "111111";
            when "0110110001110" => rgb <= "111111";
            when "0110110001111" => rgb <= "111111";
            when "0110110010000" => rgb <= "111111";
            when "0110110010001" => rgb <= "111111";
            when "0110110010010" => rgb <= "111111";
            when "0110110010011" => rgb <= "111111";
            when "0110110010100" => rgb <= "111111";
            when "0110110010101" => rgb <= "111111";
            when "0110110010110" => rgb <= "111111";
            when "0110110010111" => rgb <= "111111";
            when "0110110011000" => rgb <= "111111";
            when "0110110011001" => rgb <= "111111";
            when "0110110011010" => rgb <= "111111";
            when "0110110011011" => rgb <= "111111";
            when "0110110011100" => rgb <= "111111";
            when "0110110011101" => rgb <= "111111";
            when "0110110011110" => rgb <= "111111";
            when "0110110011111" => rgb <= "111111";
            when "0110110100000" => rgb <= "111111";
            when "0110110100001" => rgb <= "010101";
            when "0110110100010" => rgb <= "100001";
            when "0110110100011" => rgb <= "100001";
            when "0110110100100" => rgb <= "100001";
            when "0110110100101" => rgb <= "100001";
            when "0110110100110" => rgb <= "100001";
            when "0110110100111" => rgb <= "100001";
            when "0110111000000" => rgb <= "100001";
            when "0110111000001" => rgb <= "100001";
            when "0110111000010" => rgb <= "100001";
            when "0110111000011" => rgb <= "100001";
            when "0110111000100" => rgb <= "100001";
            when "0110111000101" => rgb <= "100001";
            when "0110111000110" => rgb <= "100001";
            when "0110111000111" => rgb <= "010101";
            when "0110111001000" => rgb <= "101010";
            when "0110111001001" => rgb <= "101010";
            when "0110111001010" => rgb <= "101010";
            when "0110111001011" => rgb <= "111111";
            when "0110111001100" => rgb <= "111111";
            when "0110111001101" => rgb <= "111111";
            when "0110111001110" => rgb <= "111111";
            when "0110111001111" => rgb <= "111111";
            when "0110111010000" => rgb <= "111111";
            when "0110111010001" => rgb <= "111111";
            when "0110111010010" => rgb <= "111111";
            when "0110111010011" => rgb <= "111111";
            when "0110111010100" => rgb <= "111111";
            when "0110111010101" => rgb <= "111111";
            when "0110111010110" => rgb <= "111111";
            when "0110111010111" => rgb <= "111111";
            when "0110111011000" => rgb <= "111111";
            when "0110111011001" => rgb <= "111111";
            when "0110111011010" => rgb <= "111111";
            when "0110111011011" => rgb <= "111111";
            when "0110111011100" => rgb <= "111111";
            when "0110111011101" => rgb <= "111111";
            when "0110111011110" => rgb <= "111111";
            when "0110111011111" => rgb <= "111111";
            when "0110111100000" => rgb <= "111111";
            when "0110111100001" => rgb <= "010101";
            when "0110111100010" => rgb <= "100001";
            when "0110111100011" => rgb <= "100001";
            when "0110111100100" => rgb <= "100001";
            when "0110111100101" => rgb <= "100001";
            when "0110111100110" => rgb <= "100001";
            when "0110111100111" => rgb <= "100001";
            when "0111000000000" => rgb <= "100001";
            when "0111000000001" => rgb <= "100001";
            when "0111000000010" => rgb <= "100001";
            when "0111000000011" => rgb <= "100001";
            when "0111000000100" => rgb <= "100001";
            when "0111000000101" => rgb <= "100001";
            when "0111000000110" => rgb <= "100001";
            when "0111000000111" => rgb <= "010101";
            when "0111000001000" => rgb <= "101010";
            when "0111000001001" => rgb <= "101010";
            when "0111000001010" => rgb <= "111111";
            when "0111000001011" => rgb <= "111111";
            when "0111000001100" => rgb <= "111111";
            when "0111000001101" => rgb <= "111111";
            when "0111000001110" => rgb <= "111111";
            when "0111000001111" => rgb <= "111111";
            when "0111000010000" => rgb <= "111111";
            when "0111000010001" => rgb <= "111111";
            when "0111000010010" => rgb <= "111111";
            when "0111000010011" => rgb <= "111111";
            when "0111000010100" => rgb <= "111111";
            when "0111000010101" => rgb <= "111111";
            when "0111000010110" => rgb <= "111111";
            when "0111000010111" => rgb <= "111111";
            when "0111000011000" => rgb <= "111111";
            when "0111000011001" => rgb <= "111111";
            when "0111000011010" => rgb <= "111111";
            when "0111000011011" => rgb <= "111111";
            when "0111000011100" => rgb <= "111111";
            when "0111000011101" => rgb <= "111111";
            when "0111000011110" => rgb <= "111111";
            when "0111000011111" => rgb <= "111111";
            when "0111000100000" => rgb <= "111111";
            when "0111000100001" => rgb <= "010101";
            when "0111000100010" => rgb <= "100001";
            when "0111000100011" => rgb <= "100001";
            when "0111000100100" => rgb <= "100001";
            when "0111000100101" => rgb <= "100001";
            when "0111000100110" => rgb <= "100001";
            when "0111000100111" => rgb <= "100001";
            when "0111001000000" => rgb <= "100001";
            when "0111001000001" => rgb <= "100001";
            when "0111001000010" => rgb <= "100001";
            when "0111001000011" => rgb <= "100001";
            when "0111001000100" => rgb <= "100001";
            when "0111001000101" => rgb <= "100001";
            when "0111001000110" => rgb <= "100001";
            when "0111001000111" => rgb <= "010101";
            when "0111001001000" => rgb <= "101010";
            when "0111001001001" => rgb <= "101010";
            when "0111001001010" => rgb <= "111111";
            when "0111001001011" => rgb <= "111111";
            when "0111001001100" => rgb <= "111111";
            when "0111001001101" => rgb <= "111111";
            when "0111001001110" => rgb <= "111111";
            when "0111001001111" => rgb <= "111111";
            when "0111001010000" => rgb <= "111111";
            when "0111001010001" => rgb <= "111111";
            when "0111001010010" => rgb <= "111111";
            when "0111001010011" => rgb <= "111111";
            when "0111001010100" => rgb <= "111111";
            when "0111001010101" => rgb <= "111111";
            when "0111001010110" => rgb <= "111111";
            when "0111001010111" => rgb <= "111111";
            when "0111001011000" => rgb <= "111111";
            when "0111001011001" => rgb <= "111111";
            when "0111001011010" => rgb <= "111111";
            when "0111001011011" => rgb <= "111111";
            when "0111001011100" => rgb <= "111111";
            when "0111001011101" => rgb <= "111111";
            when "0111001011110" => rgb <= "111111";
            when "0111001011111" => rgb <= "111111";
            when "0111001100000" => rgb <= "111111";
            when "0111001100001" => rgb <= "111111";
            when "0111001100010" => rgb <= "010101";
            when "0111001100011" => rgb <= "100001";
            when "0111001100100" => rgb <= "100001";
            when "0111001100101" => rgb <= "100001";
            when "0111001100110" => rgb <= "100001";
            when "0111001100111" => rgb <= "100001";
            when "0111010000000" => rgb <= "100001";
            when "0111010000001" => rgb <= "100001";
            when "0111010000010" => rgb <= "100001";
            when "0111010000011" => rgb <= "100001";
            when "0111010000100" => rgb <= "100001";
            when "0111010000101" => rgb <= "100001";
            when "0111010000110" => rgb <= "100001";
            when "0111010000111" => rgb <= "010101";
            when "0111010001000" => rgb <= "101010";
            when "0111010001001" => rgb <= "101010";
            when "0111010001010" => rgb <= "111111";
            when "0111010001011" => rgb <= "111111";
            when "0111010001100" => rgb <= "111111";
            when "0111010001101" => rgb <= "111111";
            when "0111010001110" => rgb <= "111111";
            when "0111010001111" => rgb <= "111111";
            when "0111010010000" => rgb <= "111111";
            when "0111010010001" => rgb <= "111111";
            when "0111010010010" => rgb <= "111111";
            when "0111010010011" => rgb <= "111111";
            when "0111010010100" => rgb <= "111111";
            when "0111010010101" => rgb <= "111111";
            when "0111010010110" => rgb <= "111111";
            when "0111010010111" => rgb <= "111111";
            when "0111010011000" => rgb <= "111111";
            when "0111010011001" => rgb <= "111111";
            when "0111010011010" => rgb <= "111111";
            when "0111010011011" => rgb <= "111111";
            when "0111010011100" => rgb <= "111111";
            when "0111010011101" => rgb <= "111111";
            when "0111010011110" => rgb <= "111111";
            when "0111010011111" => rgb <= "111111";
            when "0111010100000" => rgb <= "111111";
            when "0111010100001" => rgb <= "111111";
            when "0111010100010" => rgb <= "010101";
            when "0111010100011" => rgb <= "100001";
            when "0111010100100" => rgb <= "100001";
            when "0111010100101" => rgb <= "100001";
            when "0111010100110" => rgb <= "100001";
            when "0111010100111" => rgb <= "100001";
            when "0111011000000" => rgb <= "100001";
            when "0111011000001" => rgb <= "100001";
            when "0111011000010" => rgb <= "100001";
            when "0111011000011" => rgb <= "100001";
            when "0111011000100" => rgb <= "100001";
            when "0111011000101" => rgb <= "100001";
            when "0111011000110" => rgb <= "100001";
            when "0111011000111" => rgb <= "010101";
            when "0111011001000" => rgb <= "101010";
            when "0111011001001" => rgb <= "101010";
            when "0111011001010" => rgb <= "111111";
            when "0111011001011" => rgb <= "111111";
            when "0111011001100" => rgb <= "111111";
            when "0111011001101" => rgb <= "111111";
            when "0111011001110" => rgb <= "111111";
            when "0111011001111" => rgb <= "111111";
            when "0111011010000" => rgb <= "111111";
            when "0111011010001" => rgb <= "111111";
            when "0111011010010" => rgb <= "111111";
            when "0111011010011" => rgb <= "111111";
            when "0111011010100" => rgb <= "111111";
            when "0111011010101" => rgb <= "111111";
            when "0111011010110" => rgb <= "111111";
            when "0111011010111" => rgb <= "111111";
            when "0111011011000" => rgb <= "111111";
            when "0111011011001" => rgb <= "111111";
            when "0111011011010" => rgb <= "111111";
            when "0111011011011" => rgb <= "111111";
            when "0111011011100" => rgb <= "111111";
            when "0111011011101" => rgb <= "111111";
            when "0111011011110" => rgb <= "111111";
            when "0111011011111" => rgb <= "111111";
            when "0111011100000" => rgb <= "111111";
            when "0111011100001" => rgb <= "111111";
            when "0111011100010" => rgb <= "010101";
            when "0111011100011" => rgb <= "100001";
            when "0111011100100" => rgb <= "100001";
            when "0111011100101" => rgb <= "100001";
            when "0111011100110" => rgb <= "100001";
            when "0111011100111" => rgb <= "100001";
            when "0111100000000" => rgb <= "100001";
            when "0111100000001" => rgb <= "100001";
            when "0111100000010" => rgb <= "100001";
            when "0111100000011" => rgb <= "100001";
            when "0111100000100" => rgb <= "100001";
            when "0111100000101" => rgb <= "100001";
            when "0111100000110" => rgb <= "100001";
            when "0111100000111" => rgb <= "010101";
            when "0111100001000" => rgb <= "101010";
            when "0111100001001" => rgb <= "101010";
            when "0111100001010" => rgb <= "111111";
            when "0111100001011" => rgb <= "111111";
            when "0111100001100" => rgb <= "111111";
            when "0111100001101" => rgb <= "111111";
            when "0111100001110" => rgb <= "111111";
            when "0111100001111" => rgb <= "111111";
            when "0111100010000" => rgb <= "111111";
            when "0111100010001" => rgb <= "111111";
            when "0111100010010" => rgb <= "111111";
            when "0111100010011" => rgb <= "111111";
            when "0111100010100" => rgb <= "111111";
            when "0111100010101" => rgb <= "111111";
            when "0111100010110" => rgb <= "111111";
            when "0111100010111" => rgb <= "111111";
            when "0111100011000" => rgb <= "111111";
            when "0111100011001" => rgb <= "111111";
            when "0111100011010" => rgb <= "111111";
            when "0111100011011" => rgb <= "111111";
            when "0111100011100" => rgb <= "111111";
            when "0111100011101" => rgb <= "111111";
            when "0111100011110" => rgb <= "111111";
            when "0111100011111" => rgb <= "111111";
            when "0111100100000" => rgb <= "111111";
            when "0111100100001" => rgb <= "111111";
            when "0111100100010" => rgb <= "010101";
            when "0111100100011" => rgb <= "100001";
            when "0111100100100" => rgb <= "100001";
            when "0111100100101" => rgb <= "100001";
            when "0111100100110" => rgb <= "100001";
            when "0111100100111" => rgb <= "100001";
            when "0111101000000" => rgb <= "100001";
            when "0111101000001" => rgb <= "100001";
            when "0111101000010" => rgb <= "100001";
            when "0111101000011" => rgb <= "100001";
            when "0111101000100" => rgb <= "100001";
            when "0111101000101" => rgb <= "100001";
            when "0111101000110" => rgb <= "100001";
            when "0111101000111" => rgb <= "010101";
            when "0111101001000" => rgb <= "101010";
            when "0111101001001" => rgb <= "101010";
            when "0111101001010" => rgb <= "111111";
            when "0111101001011" => rgb <= "111111";
            when "0111101001100" => rgb <= "111111";
            when "0111101001101" => rgb <= "111111";
            when "0111101001110" => rgb <= "111111";
            when "0111101001111" => rgb <= "111111";
            when "0111101010000" => rgb <= "111111";
            when "0111101010001" => rgb <= "111111";
            when "0111101010010" => rgb <= "111111";
            when "0111101010011" => rgb <= "111111";
            when "0111101010100" => rgb <= "111111";
            when "0111101010101" => rgb <= "111111";
            when "0111101010110" => rgb <= "111111";
            when "0111101010111" => rgb <= "111111";
            when "0111101011000" => rgb <= "111111";
            when "0111101011001" => rgb <= "111111";
            when "0111101011010" => rgb <= "111111";
            when "0111101011011" => rgb <= "111111";
            when "0111101011100" => rgb <= "111111";
            when "0111101011101" => rgb <= "111111";
            when "0111101011110" => rgb <= "111111";
            when "0111101011111" => rgb <= "111111";
            when "0111101100000" => rgb <= "111111";
            when "0111101100001" => rgb <= "111111";
            when "0111101100010" => rgb <= "010101";
            when "0111101100011" => rgb <= "100001";
            when "0111101100100" => rgb <= "100001";
            when "0111101100101" => rgb <= "100001";
            when "0111101100110" => rgb <= "100001";
            when "0111101100111" => rgb <= "100001";
            when "0111110000000" => rgb <= "100001";
            when "0111110000001" => rgb <= "100001";
            when "0111110000010" => rgb <= "100001";
            when "0111110000011" => rgb <= "100001";
            when "0111110000100" => rgb <= "100001";
            when "0111110000101" => rgb <= "100001";
            when "0111110000110" => rgb <= "010101";
            when "0111110000111" => rgb <= "101010";
            when "0111110001000" => rgb <= "101010";
            when "0111110001001" => rgb <= "111111";
            when "0111110001010" => rgb <= "111111";
            when "0111110001011" => rgb <= "111111";
            when "0111110001100" => rgb <= "111111";
            when "0111110001101" => rgb <= "111111";
            when "0111110001110" => rgb <= "111111";
            when "0111110001111" => rgb <= "111111";
            when "0111110010000" => rgb <= "111111";
            when "0111110010001" => rgb <= "111111";
            when "0111110010010" => rgb <= "111111";
            when "0111110010011" => rgb <= "111111";
            when "0111110010100" => rgb <= "111111";
            when "0111110010101" => rgb <= "111111";
            when "0111110010110" => rgb <= "111111";
            when "0111110010111" => rgb <= "111111";
            when "0111110011000" => rgb <= "111111";
            when "0111110011001" => rgb <= "111111";
            when "0111110011010" => rgb <= "111111";
            when "0111110011011" => rgb <= "111111";
            when "0111110011100" => rgb <= "111111";
            when "0111110011101" => rgb <= "111111";
            when "0111110011110" => rgb <= "111111";
            when "0111110011111" => rgb <= "111111";
            when "0111110100000" => rgb <= "111111";
            when "0111110100001" => rgb <= "111111";
            when "0111110100010" => rgb <= "010101";
            when "0111110100011" => rgb <= "100001";
            when "0111110100100" => rgb <= "100001";
            when "0111110100101" => rgb <= "100001";
            when "0111110100110" => rgb <= "100001";
            when "0111110100111" => rgb <= "100001";
            when "0111111000000" => rgb <= "100001";
            when "0111111000001" => rgb <= "100001";
            when "0111111000010" => rgb <= "100001";
            when "0111111000011" => rgb <= "100001";
            when "0111111000100" => rgb <= "100001";
            when "0111111000101" => rgb <= "100001";
            when "0111111000110" => rgb <= "010101";
            when "0111111000111" => rgb <= "101010";
            when "0111111001000" => rgb <= "101010";
            when "0111111001001" => rgb <= "111111";
            when "0111111001010" => rgb <= "111111";
            when "0111111001011" => rgb <= "111111";
            when "0111111001100" => rgb <= "111111";
            when "0111111001101" => rgb <= "111111";
            when "0111111001110" => rgb <= "111111";
            when "0111111001111" => rgb <= "111111";
            when "0111111010000" => rgb <= "111111";
            when "0111111010001" => rgb <= "111111";
            when "0111111010010" => rgb <= "111111";
            when "0111111010011" => rgb <= "111111";
            when "0111111010100" => rgb <= "111111";
            when "0111111010101" => rgb <= "111111";
            when "0111111010110" => rgb <= "111111";
            when "0111111010111" => rgb <= "111111";
            when "0111111011000" => rgb <= "111111";
            when "0111111011001" => rgb <= "111111";
            when "0111111011010" => rgb <= "111111";
            when "0111111011011" => rgb <= "111111";
            when "0111111011100" => rgb <= "111111";
            when "0111111011101" => rgb <= "111111";
            when "0111111011110" => rgb <= "111111";
            when "0111111011111" => rgb <= "111111";
            when "0111111100000" => rgb <= "111111";
            when "0111111100001" => rgb <= "111111";
            when "0111111100010" => rgb <= "010101";
            when "0111111100011" => rgb <= "100001";
            when "0111111100100" => rgb <= "100001";
            when "0111111100101" => rgb <= "100001";
            when "0111111100110" => rgb <= "100001";
            when "0111111100111" => rgb <= "100001";
            when "1000000000000" => rgb <= "100001";
            when "1000000000001" => rgb <= "100001";
            when "1000000000010" => rgb <= "100001";
            when "1000000000011" => rgb <= "100001";
            when "1000000000100" => rgb <= "100001";
            when "1000000000101" => rgb <= "100001";
            when "1000000000110" => rgb <= "010101";
            when "1000000000111" => rgb <= "101010";
            when "1000000001000" => rgb <= "101010";
            when "1000000001001" => rgb <= "111111";
            when "1000000001010" => rgb <= "111111";
            when "1000000001011" => rgb <= "111111";
            when "1000000001100" => rgb <= "111111";
            when "1000000001101" => rgb <= "111111";
            when "1000000001110" => rgb <= "111111";
            when "1000000001111" => rgb <= "111111";
            when "1000000010000" => rgb <= "111111";
            when "1000000010001" => rgb <= "111111";
            when "1000000010010" => rgb <= "111111";
            when "1000000010011" => rgb <= "111111";
            when "1000000010100" => rgb <= "111111";
            when "1000000010101" => rgb <= "111111";
            when "1000000010110" => rgb <= "111111";
            when "1000000010111" => rgb <= "111111";
            when "1000000011000" => rgb <= "111111";
            when "1000000011001" => rgb <= "111111";
            when "1000000011010" => rgb <= "111111";
            when "1000000011011" => rgb <= "111111";
            when "1000000011100" => rgb <= "111111";
            when "1000000011101" => rgb <= "111111";
            when "1000000011110" => rgb <= "111111";
            when "1000000011111" => rgb <= "111111";
            when "1000000100000" => rgb <= "111111";
            when "1000000100001" => rgb <= "111111";
            when "1000000100010" => rgb <= "010101";
            when "1000000100011" => rgb <= "100001";
            when "1000000100100" => rgb <= "100001";
            when "1000000100101" => rgb <= "100001";
            when "1000000100110" => rgb <= "100001";
            when "1000000100111" => rgb <= "100001";
            when "1000001000000" => rgb <= "100001";
            when "1000001000001" => rgb <= "100001";
            when "1000001000010" => rgb <= "100001";
            when "1000001000011" => rgb <= "100001";
            when "1000001000100" => rgb <= "100001";
            when "1000001000101" => rgb <= "100001";
            when "1000001000110" => rgb <= "010101";
            when "1000001000111" => rgb <= "101010";
            when "1000001001000" => rgb <= "101010";
            when "1000001001001" => rgb <= "111111";
            when "1000001001010" => rgb <= "111111";
            when "1000001001011" => rgb <= "111111";
            when "1000001001100" => rgb <= "111111";
            when "1000001001101" => rgb <= "111111";
            when "1000001001110" => rgb <= "111111";
            when "1000001001111" => rgb <= "111111";
            when "1000001010000" => rgb <= "111111";
            when "1000001010001" => rgb <= "111111";
            when "1000001010010" => rgb <= "111111";
            when "1000001010011" => rgb <= "111111";
            when "1000001010100" => rgb <= "111111";
            when "1000001010101" => rgb <= "111111";
            when "1000001010110" => rgb <= "111111";
            when "1000001010111" => rgb <= "111111";
            when "1000001011000" => rgb <= "111111";
            when "1000001011001" => rgb <= "111111";
            when "1000001011010" => rgb <= "111111";
            when "1000001011011" => rgb <= "111111";
            when "1000001011100" => rgb <= "111111";
            when "1000001011101" => rgb <= "111111";
            when "1000001011110" => rgb <= "111111";
            when "1000001011111" => rgb <= "111111";
            when "1000001100000" => rgb <= "111111";
            when "1000001100001" => rgb <= "111111";
            when "1000001100010" => rgb <= "010101";
            when "1000001100011" => rgb <= "100001";
            when "1000001100100" => rgb <= "100001";
            when "1000001100101" => rgb <= "100001";
            when "1000001100110" => rgb <= "100001";
            when "1000001100111" => rgb <= "100001";
            when "1000010000000" => rgb <= "100001";
            when "1000010000001" => rgb <= "100001";
            when "1000010000010" => rgb <= "100001";
            when "1000010000011" => rgb <= "100001";
            when "1000010000100" => rgb <= "100001";
            when "1000010000101" => rgb <= "100001";
            when "1000010000110" => rgb <= "010101";
            when "1000010000111" => rgb <= "101010";
            when "1000010001000" => rgb <= "101010";
            when "1000010001001" => rgb <= "111111";
            when "1000010001010" => rgb <= "111111";
            when "1000010001011" => rgb <= "111111";
            when "1000010001100" => rgb <= "111111";
            when "1000010001101" => rgb <= "111111";
            when "1000010001110" => rgb <= "111111";
            when "1000010001111" => rgb <= "111111";
            when "1000010010000" => rgb <= "111111";
            when "1000010010001" => rgb <= "111111";
            when "1000010010010" => rgb <= "111111";
            when "1000010010011" => rgb <= "111111";
            when "1000010010100" => rgb <= "111111";
            when "1000010010101" => rgb <= "111111";
            when "1000010010110" => rgb <= "111111";
            when "1000010010111" => rgb <= "111111";
            when "1000010011000" => rgb <= "111111";
            when "1000010011001" => rgb <= "111111";
            when "1000010011010" => rgb <= "111111";
            when "1000010011011" => rgb <= "111111";
            when "1000010011100" => rgb <= "111111";
            when "1000010011101" => rgb <= "111111";
            when "1000010011110" => rgb <= "111111";
            when "1000010011111" => rgb <= "111111";
            when "1000010100000" => rgb <= "111111";
            when "1000010100001" => rgb <= "111111";
            when "1000010100010" => rgb <= "010101";
            when "1000010100011" => rgb <= "100001";
            when "1000010100100" => rgb <= "100001";
            when "1000010100101" => rgb <= "100001";
            when "1000010100110" => rgb <= "100001";
            when "1000010100111" => rgb <= "100001";
            when "1000011000000" => rgb <= "100001";
            when "1000011000001" => rgb <= "100001";
            when "1000011000010" => rgb <= "100001";
            when "1000011000011" => rgb <= "100001";
            when "1000011000100" => rgb <= "100001";
            when "1000011000101" => rgb <= "100001";
            when "1000011000110" => rgb <= "010101";
            when "1000011000111" => rgb <= "101010";
            when "1000011001000" => rgb <= "101010";
            when "1000011001001" => rgb <= "111111";
            when "1000011001010" => rgb <= "111111";
            when "1000011001011" => rgb <= "111111";
            when "1000011001100" => rgb <= "111111";
            when "1000011001101" => rgb <= "111111";
            when "1000011001110" => rgb <= "111111";
            when "1000011001111" => rgb <= "111111";
            when "1000011010000" => rgb <= "111111";
            when "1000011010001" => rgb <= "111111";
            when "1000011010010" => rgb <= "111111";
            when "1000011010011" => rgb <= "111111";
            when "1000011010100" => rgb <= "111111";
            when "1000011010101" => rgb <= "111111";
            when "1000011010110" => rgb <= "111111";
            when "1000011010111" => rgb <= "111111";
            when "1000011011000" => rgb <= "111111";
            when "1000011011001" => rgb <= "111111";
            when "1000011011010" => rgb <= "111111";
            when "1000011011011" => rgb <= "111111";
            when "1000011011100" => rgb <= "111111";
            when "1000011011101" => rgb <= "111111";
            when "1000011011110" => rgb <= "111111";
            when "1000011011111" => rgb <= "111111";
            when "1000011100000" => rgb <= "111111";
            when "1000011100001" => rgb <= "111111";
            when "1000011100010" => rgb <= "010101";
            when "1000011100011" => rgb <= "100001";
            when "1000011100100" => rgb <= "100001";
            when "1000011100101" => rgb <= "100001";
            when "1000011100110" => rgb <= "100001";
            when "1000011100111" => rgb <= "100001";
            when "1000100000000" => rgb <= "100001";
            when "1000100000001" => rgb <= "100001";
            when "1000100000010" => rgb <= "100001";
            when "1000100000011" => rgb <= "100001";
            when "1000100000100" => rgb <= "100001";
            when "1000100000101" => rgb <= "100001";
            when "1000100000110" => rgb <= "010101";
            when "1000100000111" => rgb <= "101010";
            when "1000100001000" => rgb <= "101010";
            when "1000100001001" => rgb <= "111111";
            when "1000100001010" => rgb <= "111111";
            when "1000100001011" => rgb <= "111111";
            when "1000100001100" => rgb <= "111111";
            when "1000100001101" => rgb <= "111111";
            when "1000100001110" => rgb <= "111111";
            when "1000100001111" => rgb <= "111111";
            when "1000100010000" => rgb <= "111111";
            when "1000100010001" => rgb <= "111111";
            when "1000100010010" => rgb <= "111111";
            when "1000100010011" => rgb <= "111111";
            when "1000100010100" => rgb <= "111111";
            when "1000100010101" => rgb <= "111111";
            when "1000100010110" => rgb <= "111111";
            when "1000100010111" => rgb <= "111111";
            when "1000100011000" => rgb <= "111111";
            when "1000100011001" => rgb <= "111111";
            when "1000100011010" => rgb <= "111111";
            when "1000100011011" => rgb <= "111111";
            when "1000100011100" => rgb <= "111111";
            when "1000100011101" => rgb <= "111111";
            when "1000100011110" => rgb <= "111111";
            when "1000100011111" => rgb <= "111111";
            when "1000100100000" => rgb <= "111111";
            when "1000100100001" => rgb <= "111111";
            when "1000100100010" => rgb <= "010101";
            when "1000100100011" => rgb <= "100001";
            when "1000100100100" => rgb <= "100001";
            when "1000100100101" => rgb <= "100001";
            when "1000100100110" => rgb <= "100001";
            when "1000100100111" => rgb <= "100001";
            when "1000101000000" => rgb <= "100001";
            when "1000101000001" => rgb <= "100001";
            when "1000101000010" => rgb <= "100001";
            when "1000101000011" => rgb <= "100001";
            when "1000101000100" => rgb <= "100001";
            when "1000101000101" => rgb <= "100001";
            when "1000101000110" => rgb <= "010101";
            when "1000101000111" => rgb <= "101010";
            when "1000101001000" => rgb <= "101010";
            when "1000101001001" => rgb <= "111111";
            when "1000101001010" => rgb <= "111111";
            when "1000101001011" => rgb <= "111111";
            when "1000101001100" => rgb <= "111111";
            when "1000101001101" => rgb <= "111111";
            when "1000101001110" => rgb <= "111111";
            when "1000101001111" => rgb <= "111111";
            when "1000101010000" => rgb <= "111111";
            when "1000101010001" => rgb <= "111111";
            when "1000101010010" => rgb <= "111111";
            when "1000101010011" => rgb <= "111111";
            when "1000101010100" => rgb <= "111111";
            when "1000101010101" => rgb <= "111111";
            when "1000101010110" => rgb <= "111111";
            when "1000101010111" => rgb <= "111111";
            when "1000101011000" => rgb <= "111111";
            when "1000101011001" => rgb <= "111111";
            when "1000101011010" => rgb <= "111111";
            when "1000101011011" => rgb <= "111111";
            when "1000101011100" => rgb <= "111111";
            when "1000101011101" => rgb <= "111111";
            when "1000101011110" => rgb <= "111111";
            when "1000101011111" => rgb <= "111111";
            when "1000101100000" => rgb <= "111111";
            when "1000101100001" => rgb <= "111111";
            when "1000101100010" => rgb <= "010101";
            when "1000101100011" => rgb <= "100001";
            when "1000101100100" => rgb <= "100001";
            when "1000101100101" => rgb <= "100001";
            when "1000101100110" => rgb <= "100001";
            when "1000101100111" => rgb <= "100001";
            when "1000110000000" => rgb <= "100001";
            when "1000110000001" => rgb <= "100001";
            when "1000110000010" => rgb <= "100001";
            when "1000110000011" => rgb <= "100001";
            when "1000110000100" => rgb <= "100001";
            when "1000110000101" => rgb <= "100001";
            when "1000110000110" => rgb <= "100001";
            when "1000110000111" => rgb <= "010101";
            when "1000110001000" => rgb <= "101010";
            when "1000110001001" => rgb <= "101010";
            when "1000110001010" => rgb <= "111111";
            when "1000110001011" => rgb <= "111111";
            when "1000110001100" => rgb <= "111111";
            when "1000110001101" => rgb <= "111111";
            when "1000110001110" => rgb <= "111111";
            when "1000110001111" => rgb <= "111111";
            when "1000110010000" => rgb <= "111111";
            when "1000110010001" => rgb <= "111111";
            when "1000110010010" => rgb <= "111111";
            when "1000110010011" => rgb <= "111111";
            when "1000110010100" => rgb <= "111111";
            when "1000110010101" => rgb <= "111111";
            when "1000110010110" => rgb <= "111111";
            when "1000110010111" => rgb <= "111111";
            when "1000110011000" => rgb <= "111111";
            when "1000110011001" => rgb <= "111111";
            when "1000110011010" => rgb <= "111111";
            when "1000110011011" => rgb <= "111111";
            when "1000110011100" => rgb <= "111111";
            when "1000110011101" => rgb <= "111111";
            when "1000110011110" => rgb <= "111111";
            when "1000110011111" => rgb <= "111111";
            when "1000110100000" => rgb <= "111111";
            when "1000110100001" => rgb <= "111111";
            when "1000110100010" => rgb <= "010101";
            when "1000110100011" => rgb <= "100001";
            when "1000110100100" => rgb <= "100001";
            when "1000110100101" => rgb <= "100001";
            when "1000110100110" => rgb <= "100001";
            when "1000110100111" => rgb <= "100001";
            when "1000111000000" => rgb <= "100001";
            when "1000111000001" => rgb <= "100001";
            when "1000111000010" => rgb <= "100001";
            when "1000111000011" => rgb <= "100001";
            when "1000111000100" => rgb <= "100001";
            when "1000111000101" => rgb <= "100001";
            when "1000111000110" => rgb <= "100001";
            when "1000111000111" => rgb <= "100001";
            when "1000111001000" => rgb <= "010101";
            when "1000111001001" => rgb <= "101010";
            when "1000111001010" => rgb <= "101010";
            when "1000111001011" => rgb <= "111111";
            when "1000111001100" => rgb <= "111111";
            when "1000111001101" => rgb <= "111111";
            when "1000111001110" => rgb <= "111111";
            when "1000111001111" => rgb <= "111111";
            when "1000111010000" => rgb <= "111111";
            when "1000111010001" => rgb <= "111111";
            when "1000111010010" => rgb <= "111111";
            when "1000111010011" => rgb <= "111111";
            when "1000111010100" => rgb <= "111111";
            when "1000111010101" => rgb <= "111111";
            when "1000111010110" => rgb <= "111111";
            when "1000111010111" => rgb <= "111111";
            when "1000111011000" => rgb <= "111111";
            when "1000111011001" => rgb <= "111111";
            when "1000111011010" => rgb <= "111111";
            when "1000111011011" => rgb <= "111111";
            when "1000111011100" => rgb <= "111111";
            when "1000111011101" => rgb <= "111111";
            when "1000111011110" => rgb <= "111111";
            when "1000111011111" => rgb <= "111111";
            when "1000111100000" => rgb <= "111111";
            when "1000111100001" => rgb <= "010101";
            when "1000111100010" => rgb <= "100001";
            when "1000111100011" => rgb <= "100001";
            when "1000111100100" => rgb <= "100001";
            when "1000111100101" => rgb <= "100001";
            when "1000111100110" => rgb <= "100001";
            when "1000111100111" => rgb <= "100001";
            when "1001000000000" => rgb <= "100001";
            when "1001000000001" => rgb <= "100001";
            when "1001000000010" => rgb <= "100001";
            when "1001000000011" => rgb <= "100001";
            when "1001000000100" => rgb <= "100001";
            when "1001000000101" => rgb <= "100001";
            when "1001000000110" => rgb <= "100001";
            when "1001000000111" => rgb <= "100001";
            when "1001000001000" => rgb <= "100001";
            when "1001000001001" => rgb <= "010101";
            when "1001000001010" => rgb <= "101010";
            when "1001000001011" => rgb <= "101010";
            when "1001000001100" => rgb <= "111111";
            when "1001000001101" => rgb <= "111111";
            when "1001000001110" => rgb <= "111111";
            when "1001000001111" => rgb <= "111111";
            when "1001000010000" => rgb <= "111111";
            when "1001000010001" => rgb <= "111111";
            when "1001000010010" => rgb <= "111111";
            when "1001000010011" => rgb <= "111111";
            when "1001000010100" => rgb <= "111111";
            when "1001000010101" => rgb <= "111111";
            when "1001000010110" => rgb <= "111111";
            when "1001000010111" => rgb <= "111111";
            when "1001000011000" => rgb <= "111111";
            when "1001000011001" => rgb <= "111111";
            when "1001000011010" => rgb <= "111111";
            when "1001000011011" => rgb <= "111111";
            when "1001000011100" => rgb <= "111111";
            when "1001000011101" => rgb <= "111111";
            when "1001000011110" => rgb <= "111111";
            when "1001000011111" => rgb <= "111111";
            when "1001000100000" => rgb <= "010101";
            when "1001000100001" => rgb <= "100001";
            when "1001000100010" => rgb <= "100001";
            when "1001000100011" => rgb <= "100001";
            when "1001000100100" => rgb <= "100001";
            when "1001000100101" => rgb <= "100001";
            when "1001000100110" => rgb <= "100001";
            when "1001000100111" => rgb <= "100001";
            when "1001001000000" => rgb <= "100001";
            when "1001001000001" => rgb <= "100001";
            when "1001001000010" => rgb <= "100001";
            when "1001001000011" => rgb <= "100001";
            when "1001001000100" => rgb <= "100001";
            when "1001001000101" => rgb <= "100001";
            when "1001001000110" => rgb <= "100001";
            when "1001001000111" => rgb <= "100001";
            when "1001001001000" => rgb <= "100001";
            when "1001001001001" => rgb <= "010101";
            when "1001001001010" => rgb <= "101010";
            when "1001001001011" => rgb <= "101010";
            when "1001001001100" => rgb <= "111111";
            when "1001001001101" => rgb <= "111111";
            when "1001001001110" => rgb <= "111111";
            when "1001001001111" => rgb <= "111111";
            when "1001001010000" => rgb <= "111111";
            when "1001001010001" => rgb <= "111111";
            when "1001001010010" => rgb <= "111111";
            when "1001001010011" => rgb <= "111111";
            when "1001001010100" => rgb <= "111111";
            when "1001001010101" => rgb <= "111111";
            when "1001001010110" => rgb <= "111111";
            when "1001001010111" => rgb <= "111111";
            when "1001001011000" => rgb <= "111111";
            when "1001001011001" => rgb <= "111111";
            when "1001001011010" => rgb <= "111111";
            when "1001001011011" => rgb <= "111111";
            when "1001001011100" => rgb <= "111111";
            when "1001001011101" => rgb <= "111111";
            when "1001001011110" => rgb <= "111111";
            when "1001001011111" => rgb <= "111111";
            when "1001001100000" => rgb <= "010101";
            when "1001001100001" => rgb <= "100001";
            when "1001001100010" => rgb <= "100001";
            when "1001001100011" => rgb <= "100001";
            when "1001001100100" => rgb <= "100001";
            when "1001001100101" => rgb <= "100001";
            when "1001001100110" => rgb <= "100001";
            when "1001001100111" => rgb <= "100001";
            when "1001010000000" => rgb <= "100001";
            when "1001010000001" => rgb <= "100001";
            when "1001010000010" => rgb <= "100001";
            when "1001010000011" => rgb <= "100001";
            when "1001010000100" => rgb <= "100001";
            when "1001010000101" => rgb <= "100001";
            when "1001010000110" => rgb <= "100001";
            when "1001010000111" => rgb <= "100001";
            when "1001010001000" => rgb <= "100001";
            when "1001010001001" => rgb <= "100001";
            when "1001010001010" => rgb <= "010101";
            when "1001010001011" => rgb <= "101010";
            when "1001010001100" => rgb <= "101010";
            when "1001010001101" => rgb <= "111111";
            when "1001010001110" => rgb <= "111111";
            when "1001010001111" => rgb <= "111111";
            when "1001010010000" => rgb <= "111111";
            when "1001010010001" => rgb <= "111111";
            when "1001010010010" => rgb <= "111111";
            when "1001010010011" => rgb <= "111111";
            when "1001010010100" => rgb <= "111111";
            when "1001010010101" => rgb <= "111111";
            when "1001010010110" => rgb <= "111111";
            when "1001010010111" => rgb <= "111111";
            when "1001010011000" => rgb <= "111111";
            when "1001010011001" => rgb <= "111111";
            when "1001010011010" => rgb <= "111111";
            when "1001010011011" => rgb <= "111111";
            when "1001010011100" => rgb <= "111111";
            when "1001010011101" => rgb <= "111111";
            when "1001010011110" => rgb <= "111111";
            when "1001010011111" => rgb <= "010101";
            when "1001010100000" => rgb <= "100001";
            when "1001010100001" => rgb <= "100001";
            when "1001010100010" => rgb <= "100001";
            when "1001010100011" => rgb <= "100001";
            when "1001010100100" => rgb <= "100001";
            when "1001010100101" => rgb <= "100001";
            when "1001010100110" => rgb <= "100001";
            when "1001010100111" => rgb <= "100001";
            when others => rgb <= "100001";
			end case;
	end if;
	end process;
	pxl <= std_logic_vector(y_cord) & std_logic_vector(x_cord);
end;