
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity p2win_rom is
	port(
		  clk : in std_logic;
		  x_cord: in unsigned(5 downto 0);
		  y_cord : in unsigned(4 downto 0); -- 0-1023
		  rgb : out std_logic_vector(5 downto 0)
	);
end p2win_rom;

architecture synth of p2win_rom is
signal totaladr : std_logic_vector(10 downto 0);
begin
   process (clk) begin
	if rising_edge(clk) then
		case totaladr is
		    when "0000000000000" => rgb <= "000000";
        when "0000000000001" => rgb <= "000000";
        when "0000000000010" => rgb <= "000000";
        when "0000000000011" => rgb <= "000000";
        when "0000000000100" => rgb <= "000000";
        when "0000000000101" => rgb <= "000000";
        when "0000000000110" => rgb <= "000000";
        when "0000000000111" => rgb <= "000000";
        when "0000000001000" => rgb <= "000000";
        when "0000000001001" => rgb <= "000000";
        when "0000000001010" => rgb <= "000000";
        when "0000000001011" => rgb <= "000000";
        when "0000000001100" => rgb <= "000000";
        when "0000000001101" => rgb <= "000000";
        when "0000000001110" => rgb <= "000000";
        when "0000000001111" => rgb <= "000000";
        when "0000000010000" => rgb <= "000000";
        when "0000000010001" => rgb <= "000000";
        when "0000000010010" => rgb <= "000000";
        when "0000000010011" => rgb <= "000000";
        when "0000000010100" => rgb <= "000000";
        when "0000000010101" => rgb <= "000000";
        when "0000000010110" => rgb <= "000000";
        when "0000000010111" => rgb <= "000000";
        when "0000000011000" => rgb <= "000000";
        when "0000000011001" => rgb <= "000000";
        when "0000000011010" => rgb <= "000000";
        when "0000000011011" => rgb <= "000000";
        when "0000000011100" => rgb <= "000000";
        when "0000000011101" => rgb <= "000000";
        when "0000000011110" => rgb <= "000000";
        when "0000000011111" => rgb <= "000000";
        when "0000000100000" => rgb <= "000000";
        when "0000000100001" => rgb <= "000000";
        when "0000000100010" => rgb <= "000000";
        when "0000000100011" => rgb <= "000000";
        when "0000000100100" => rgb <= "000000";
        when "0000000100101" => rgb <= "000000";
        when "0000000100110" => rgb <= "000000";
        when "0000000100111" => rgb <= "000000";
        when "0000001000000" => rgb <= "000000";
        when "0000001000001" => rgb <= "000000";
        when "0000001000010" => rgb <= "000000";
        when "0000001000011" => rgb <= "000000";
        when "0000001000100" => rgb <= "000000";
        when "0000001000101" => rgb <= "000000";
        when "0000001000110" => rgb <= "000000";
        when "0000001000111" => rgb <= "000000";
        when "0000001001000" => rgb <= "000000";
        when "0000001001001" => rgb <= "000000";
        when "0000001001010" => rgb <= "000000";
        when "0000001001011" => rgb <= "000000";
        when "0000001001100" => rgb <= "000000";
        when "0000001001101" => rgb <= "000000";
        when "0000001001110" => rgb <= "000000";
        when "0000001001111" => rgb <= "000000";
        when "0000001010000" => rgb <= "000000";
        when "0000001010001" => rgb <= "000000";
        when "0000001010010" => rgb <= "000000";
        when "0000001010011" => rgb <= "000000";
        when "0000001010100" => rgb <= "000000";
        when "0000001010101" => rgb <= "000000";
        when "0000001010110" => rgb <= "000000";
        when "0000001010111" => rgb <= "000000";
        when "0000001011000" => rgb <= "000000";
        when "0000001011001" => rgb <= "000000";
        when "0000001011010" => rgb <= "000000";
        when "0000001011011" => rgb <= "000000";
        when "0000001011100" => rgb <= "000000";
        when "0000001011101" => rgb <= "000000";
        when "0000001011110" => rgb <= "000000";
        when "0000001011111" => rgb <= "000000";
        when "0000001100000" => rgb <= "000000";
        when "0000001100001" => rgb <= "000000";
        when "0000001100010" => rgb <= "000000";
        when "0000001100011" => rgb <= "000000";
        when "0000001100100" => rgb <= "000000";
        when "0000001100101" => rgb <= "000000";
        when "0000001100110" => rgb <= "000000";
        when "0000001100111" => rgb <= "000000";
        when "0000010000000" => rgb <= "000000";
        when "0000010000001" => rgb <= "000000";
        when "0000010000010" => rgb <= "000000";
        when "0000010000011" => rgb <= "000000";
        when "0000010000100" => rgb <= "000000";
        when "0000010000101" => rgb <= "000000";
        when "0000010000110" => rgb <= "000000";
        when "0000010000111" => rgb <= "000000";
        when "0000010001000" => rgb <= "000000";
        when "0000010001001" => rgb <= "000000";
        when "0000010001010" => rgb <= "000000";
        when "0000010001011" => rgb <= "000000";
        when "0000010001100" => rgb <= "000000";
        when "0000010001101" => rgb <= "000000";
        when "0000010001110" => rgb <= "000000";
        when "0000010001111" => rgb <= "000000";
        when "0000010010000" => rgb <= "000000";
        when "0000010010001" => rgb <= "000000";
        when "0000010010010" => rgb <= "000000";
        when "0000010010011" => rgb <= "000000";
        when "0000010010100" => rgb <= "000000";
        when "0000010010101" => rgb <= "000000";
        when "0000010010110" => rgb <= "000000";
        when "0000010010111" => rgb <= "000000";
        when "0000010011000" => rgb <= "000000";
        when "0000010011001" => rgb <= "000000";
        when "0000010011010" => rgb <= "000000";
        when "0000010011011" => rgb <= "000000";
        when "0000010011100" => rgb <= "000000";
        when "0000010011101" => rgb <= "000000";
        when "0000010011110" => rgb <= "000000";
        when "0000010011111" => rgb <= "000000";
        when "0000010100000" => rgb <= "000000";
        when "0000010100001" => rgb <= "000000";
        when "0000010100010" => rgb <= "000000";
        when "0000010100011" => rgb <= "000000";
        when "0000010100100" => rgb <= "000000";
        when "0000010100101" => rgb <= "000000";
        when "0000010100110" => rgb <= "000000";
        when "0000010100111" => rgb <= "000000";
        when "0000011000000" => rgb <= "000000";
        when "0000011000001" => rgb <= "000000";
        when "0000011000010" => rgb <= "000000";
        when "0000011000011" => rgb <= "000000";
        when "0000011000100" => rgb <= "000000";
        when "0000011000101" => rgb <= "000000";
        when "0000011000110" => rgb <= "000000";
        when "0000011000111" => rgb <= "000000";
        when "0000011001000" => rgb <= "000000";
        when "0000011001001" => rgb <= "000000";
        when "0000011001010" => rgb <= "000000";
        when "0000011001011" => rgb <= "000000";
        when "0000011001100" => rgb <= "000000";
        when "0000011001101" => rgb <= "000000";
        when "0000011001110" => rgb <= "000000";
        when "0000011001111" => rgb <= "000000";
        when "0000011010000" => rgb <= "000000";
        when "0000011010001" => rgb <= "000000";
        when "0000011010010" => rgb <= "000000";
        when "0000011010011" => rgb <= "000000";
        when "0000011010100" => rgb <= "000000";
        when "0000011010101" => rgb <= "000000";
        when "0000011010110" => rgb <= "000000";
        when "0000011010111" => rgb <= "000000";
        when "0000011011000" => rgb <= "000000";
        when "0000011011001" => rgb <= "000000";
        when "0000011011010" => rgb <= "000000";
        when "0000011011011" => rgb <= "000000";
        when "0000011011100" => rgb <= "000000";
        when "0000011011101" => rgb <= "000000";
        when "0000011011110" => rgb <= "000000";
        when "0000011011111" => rgb <= "000000";
        when "0000011100000" => rgb <= "000000";
        when "0000011100001" => rgb <= "000000";
        when "0000011100010" => rgb <= "000000";
        when "0000011100011" => rgb <= "000000";
        when "0000011100100" => rgb <= "000000";
        when "0000011100101" => rgb <= "000000";
        when "0000011100110" => rgb <= "000000";
        when "0000011100111" => rgb <= "000000";
        when "0000100000000" => rgb <= "000000";
        when "0000100000001" => rgb <= "000000";
        when "0000100000010" => rgb <= "000000";
        when "0000100000011" => rgb <= "100000";
        when "0000100000100" => rgb <= "100000";
        when "0000100000101" => rgb <= "100000";
        when "0000100000110" => rgb <= "000000";
        when "0000100000111" => rgb <= "000000";
        when "0000100001000" => rgb <= "100000";
        when "0000100001001" => rgb <= "000000";
        when "0000100001010" => rgb <= "000000";
        when "0000100001011" => rgb <= "000000";
        when "0000100001100" => rgb <= "000000";
        when "0000100001101" => rgb <= "000000";
        when "0000100001110" => rgb <= "100000";
        when "0000100001111" => rgb <= "000000";
        when "0000100010000" => rgb <= "000000";
        when "0000100010001" => rgb <= "000000";
        when "0000100010010" => rgb <= "100000";
        when "0000100010011" => rgb <= "000000";
        when "0000100010100" => rgb <= "000000";
        when "0000100010101" => rgb <= "000000";
        when "0000100010110" => rgb <= "100000";
        when "0000100010111" => rgb <= "000000";
        when "0000100011000" => rgb <= "100000";
        when "0000100011001" => rgb <= "100000";
        when "0000100011010" => rgb <= "100000";
        when "0000100011011" => rgb <= "100000";
        when "0000100011100" => rgb <= "000000";
        when "0000100011101" => rgb <= "100000";
        when "0000100011110" => rgb <= "100000";
        when "0000100011111" => rgb <= "100000";
        when "0000100100000" => rgb <= "000000";
        when "0000100100001" => rgb <= "000000";
        when "0000100100010" => rgb <= "000000";
        when "0000100100011" => rgb <= "000000";
        when "0000100100100" => rgb <= "100000";
        when "0000100100101" => rgb <= "000000";
        when "0000100100110" => rgb <= "000000";
        when "0000100100111" => rgb <= "000000";
        when "0000101000000" => rgb <= "000000";
        when "0000101000001" => rgb <= "000000";
        when "0000101000010" => rgb <= "000000";
        when "0000101000011" => rgb <= "100000";
        when "0000101000100" => rgb <= "000000";
        when "0000101000101" => rgb <= "000000";
        when "0000101000110" => rgb <= "100000";
        when "0000101000111" => rgb <= "000000";
        when "0000101001000" => rgb <= "100000";
        when "0000101001001" => rgb <= "000000";
        when "0000101001010" => rgb <= "000000";
        when "0000101001011" => rgb <= "000000";
        when "0000101001100" => rgb <= "000000";
        when "0000101001101" => rgb <= "000000";
        when "0000101001110" => rgb <= "100000";
        when "0000101001111" => rgb <= "000000";
        when "0000101010000" => rgb <= "000000";
        when "0000101010001" => rgb <= "000000";
        when "0000101010010" => rgb <= "100000";
        when "0000101010011" => rgb <= "000000";
        when "0000101010100" => rgb <= "000000";
        when "0000101010101" => rgb <= "000000";
        when "0000101010110" => rgb <= "100000";
        when "0000101010111" => rgb <= "000000";
        when "0000101011000" => rgb <= "100000";
        when "0000101011001" => rgb <= "000000";
        when "0000101011010" => rgb <= "000000";
        when "0000101011011" => rgb <= "000000";
        when "0000101011100" => rgb <= "000000";
        when "0000101011101" => rgb <= "100000";
        when "0000101011110" => rgb <= "000000";
        when "0000101011111" => rgb <= "000000";
        when "0000101100000" => rgb <= "100000";
        when "0000101100001" => rgb <= "000000";
        when "0000101100010" => rgb <= "000000";
        when "0000101100011" => rgb <= "100000";
        when "0000101100100" => rgb <= "100000";
        when "0000101100101" => rgb <= "000000";
        when "0000101100110" => rgb <= "000000";
        when "0000101100111" => rgb <= "000000";
        when "0000110000000" => rgb <= "000000";
        when "0000110000001" => rgb <= "000000";
        when "0000110000010" => rgb <= "000000";
        when "0000110000011" => rgb <= "100000";
        when "0000110000100" => rgb <= "000000";
        when "0000110000101" => rgb <= "000000";
        when "0000110000110" => rgb <= "100000";
        when "0000110000111" => rgb <= "000000";
        when "0000110001000" => rgb <= "100000";
        when "0000110001001" => rgb <= "000000";
        when "0000110001010" => rgb <= "000000";
        when "0000110001011" => rgb <= "000000";
        when "0000110001100" => rgb <= "000000";
        when "0000110001101" => rgb <= "100000";
        when "0000110001110" => rgb <= "100000";
        when "0000110001111" => rgb <= "100000";
        when "0000110010000" => rgb <= "000000";
        when "0000110010001" => rgb <= "000000";
        when "0000110010010" => rgb <= "000000";
        when "0000110010011" => rgb <= "100000";
        when "0000110010100" => rgb <= "000000";
        when "0000110010101" => rgb <= "100000";
        when "0000110010110" => rgb <= "000000";
        when "0000110010111" => rgb <= "000000";
        when "0000110011000" => rgb <= "100000";
        when "0000110011001" => rgb <= "000000";
        when "0000110011010" => rgb <= "000000";
        when "0000110011011" => rgb <= "000000";
        when "0000110011100" => rgb <= "000000";
        when "0000110011101" => rgb <= "100000";
        when "0000110011110" => rgb <= "000000";
        when "0000110011111" => rgb <= "000000";
        when "0000110100000" => rgb <= "100000";
        when "0000110100001" => rgb <= "000000";
        when "0000110100010" => rgb <= "100000";
        when "0000110100011" => rgb <= "000000";
        when "0000110100100" => rgb <= "100000";
        when "0000110100101" => rgb <= "000000";
        when "0000110100110" => rgb <= "000000";
        when "0000110100111" => rgb <= "000000";
        when "0000111000000" => rgb <= "000000";
        when "0000111000001" => rgb <= "000000";
        when "0000111000010" => rgb <= "000000";
        when "0000111000011" => rgb <= "100000";
        when "0000111000100" => rgb <= "000000";
        when "0000111000101" => rgb <= "000000";
        when "0000111000110" => rgb <= "100000";
        when "0000111000111" => rgb <= "000000";
        when "0000111001000" => rgb <= "100000";
        when "0000111001001" => rgb <= "000000";
        when "0000111001010" => rgb <= "000000";
        when "0000111001011" => rgb <= "000000";
        when "0000111001100" => rgb <= "000000";
        when "0000111001101" => rgb <= "100000";
        when "0000111001110" => rgb <= "000000";
        when "0000111001111" => rgb <= "100000";
        when "0000111010000" => rgb <= "000000";
        when "0000111010001" => rgb <= "000000";
        when "0000111010010" => rgb <= "000000";
        when "0000111010011" => rgb <= "100000";
        when "0000111010100" => rgb <= "000000";
        when "0000111010101" => rgb <= "100000";
        when "0000111010110" => rgb <= "000000";
        when "0000111010111" => rgb <= "000000";
        when "0000111011000" => rgb <= "100000";
        when "0000111011001" => rgb <= "100000";
        when "0000111011010" => rgb <= "100000";
        when "0000111011011" => rgb <= "000000";
        when "0000111011100" => rgb <= "000000";
        when "0000111011101" => rgb <= "100000";
        when "0000111011110" => rgb <= "000000";
        when "0000111011111" => rgb <= "000000";
        when "0000111100000" => rgb <= "100000";
        when "0000111100001" => rgb <= "000000";
        when "0000111100010" => rgb <= "000000";
        when "0000111100011" => rgb <= "000000";
        when "0000111100100" => rgb <= "100000";
        when "0000111100101" => rgb <= "000000";
        when "0000111100110" => rgb <= "000000";
        when "0000111100111" => rgb <= "000000";
        when "0001000000000" => rgb <= "000000";
        when "0001000000001" => rgb <= "000000";
        when "0001000000010" => rgb <= "000000";
        when "0001000000011" => rgb <= "100000";
        when "0001000000100" => rgb <= "100000";
        when "0001000000101" => rgb <= "100000";
        when "0001000000110" => rgb <= "000000";
        when "0001000000111" => rgb <= "000000";
        when "0001000001000" => rgb <= "100000";
        when "0001000001001" => rgb <= "000000";
        when "0001000001010" => rgb <= "000000";
        when "0001000001011" => rgb <= "000000";
        when "0001000001100" => rgb <= "100000";
        when "0001000001101" => rgb <= "100000";
        when "0001000001110" => rgb <= "000000";
        when "0001000001111" => rgb <= "100000";
        when "0001000010000" => rgb <= "100000";
        when "0001000010001" => rgb <= "000000";
        when "0001000010010" => rgb <= "000000";
        when "0001000010011" => rgb <= "000000";
        when "0001000010100" => rgb <= "100000";
        when "0001000010101" => rgb <= "000000";
        when "0001000010110" => rgb <= "000000";
        when "0001000010111" => rgb <= "000000";
        when "0001000011000" => rgb <= "100000";
        when "0001000011001" => rgb <= "000000";
        when "0001000011010" => rgb <= "000000";
        when "0001000011011" => rgb <= "000000";
        when "0001000011100" => rgb <= "000000";
        when "0001000011101" => rgb <= "100000";
        when "0001000011110" => rgb <= "100000";
        when "0001000011111" => rgb <= "100000";
        when "0001000100000" => rgb <= "000000";
        when "0001000100001" => rgb <= "000000";
        when "0001000100010" => rgb <= "000000";
        when "0001000100011" => rgb <= "000000";
        when "0001000100100" => rgb <= "100000";
        when "0001000100101" => rgb <= "000000";
        when "0001000100110" => rgb <= "000000";
        when "0001000100111" => rgb <= "000000";
        when "0001001000000" => rgb <= "000000";
        when "0001001000001" => rgb <= "000000";
        when "0001001000010" => rgb <= "000000";
        when "0001001000011" => rgb <= "100000";
        when "0001001000100" => rgb <= "000000";
        when "0001001000101" => rgb <= "000000";
        when "0001001000110" => rgb <= "000000";
        when "0001001000111" => rgb <= "000000";
        when "0001001001000" => rgb <= "100000";
        when "0001001001001" => rgb <= "000000";
        when "0001001001010" => rgb <= "000000";
        when "0001001001011" => rgb <= "000000";
        when "0001001001100" => rgb <= "100000";
        when "0001001001101" => rgb <= "100000";
        when "0001001001110" => rgb <= "100000";
        when "0001001001111" => rgb <= "100000";
        when "0001001010000" => rgb <= "100000";
        when "0001001010001" => rgb <= "000000";
        when "0001001010010" => rgb <= "000000";
        when "0001001010011" => rgb <= "000000";
        when "0001001010100" => rgb <= "100000";
        when "0001001010101" => rgb <= "000000";
        when "0001001010110" => rgb <= "000000";
        when "0001001010111" => rgb <= "000000";
        when "0001001011000" => rgb <= "100000";
        when "0001001011001" => rgb <= "000000";
        when "0001001011010" => rgb <= "000000";
        when "0001001011011" => rgb <= "000000";
        when "0001001011100" => rgb <= "000000";
        when "0001001011101" => rgb <= "100000";
        when "0001001011110" => rgb <= "000000";
        when "0001001011111" => rgb <= "000000";
        when "0001001100000" => rgb <= "100000";
        when "0001001100001" => rgb <= "000000";
        when "0001001100010" => rgb <= "000000";
        when "0001001100011" => rgb <= "000000";
        when "0001001100100" => rgb <= "100000";
        when "0001001100101" => rgb <= "000000";
        when "0001001100110" => rgb <= "000000";
        when "0001001100111" => rgb <= "000000";
        when "0001010000000" => rgb <= "000000";
        when "0001010000001" => rgb <= "000000";
        when "0001010000010" => rgb <= "000000";
        when "0001010000011" => rgb <= "100000";
        when "0001010000100" => rgb <= "000000";
        when "0001010000101" => rgb <= "000000";
        when "0001010000110" => rgb <= "000000";
        when "0001010000111" => rgb <= "000000";
        when "0001010001000" => rgb <= "100000";
        when "0001010001001" => rgb <= "000000";
        when "0001010001010" => rgb <= "000000";
        when "0001010001011" => rgb <= "000000";
        when "0001010001100" => rgb <= "100000";
        when "0001010001101" => rgb <= "000000";
        when "0001010001110" => rgb <= "000000";
        when "0001010001111" => rgb <= "000000";
        when "0001010010000" => rgb <= "100000";
        when "0001010010001" => rgb <= "000000";
        when "0001010010010" => rgb <= "000000";
        when "0001010010011" => rgb <= "000000";
        when "0001010010100" => rgb <= "100000";
        when "0001010010101" => rgb <= "000000";
        when "0001010010110" => rgb <= "000000";
        when "0001010010111" => rgb <= "000000";
        when "0001010011000" => rgb <= "100000";
        when "0001010011001" => rgb <= "000000";
        when "0001010011010" => rgb <= "000000";
        when "0001010011011" => rgb <= "000000";
        when "0001010011100" => rgb <= "000000";
        when "0001010011101" => rgb <= "100000";
        when "0001010011110" => rgb <= "000000";
        when "0001010011111" => rgb <= "000000";
        when "0001010100000" => rgb <= "100000";
        when "0001010100001" => rgb <= "000000";
        when "0001010100010" => rgb <= "000000";
        when "0001010100011" => rgb <= "000000";
        when "0001010100100" => rgb <= "100000";
        when "0001010100101" => rgb <= "000000";
        when "0001010100110" => rgb <= "000000";
        when "0001010100111" => rgb <= "000000";
        when "0001011000000" => rgb <= "000000";
        when "0001011000001" => rgb <= "000000";
        when "0001011000010" => rgb <= "000000";
        when "0001011000011" => rgb <= "100000";
        when "0001011000100" => rgb <= "000000";
        when "0001011000101" => rgb <= "000000";
        when "0001011000110" => rgb <= "000000";
        when "0001011000111" => rgb <= "000000";
        when "0001011001000" => rgb <= "100000";
        when "0001011001001" => rgb <= "100000";
        when "0001011001010" => rgb <= "100000";
        when "0001011001011" => rgb <= "000000";
        when "0001011001100" => rgb <= "100000";
        when "0001011001101" => rgb <= "000000";
        when "0001011001110" => rgb <= "000000";
        when "0001011001111" => rgb <= "000000";
        when "0001011010000" => rgb <= "100000";
        when "0001011010001" => rgb <= "000000";
        when "0001011010010" => rgb <= "000000";
        when "0001011010011" => rgb <= "000000";
        when "0001011010100" => rgb <= "100000";
        when "0001011010101" => rgb <= "000000";
        when "0001011010110" => rgb <= "000000";
        when "0001011010111" => rgb <= "000000";
        when "0001011011000" => rgb <= "100000";
        when "0001011011001" => rgb <= "100000";
        when "0001011011010" => rgb <= "100000";
        when "0001011011011" => rgb <= "100000";
        when "0001011011100" => rgb <= "000000";
        when "0001011011101" => rgb <= "100000";
        when "0001011011110" => rgb <= "000000";
        when "0001011011111" => rgb <= "000000";
        when "0001011100000" => rgb <= "100000";
        when "0001011100001" => rgb <= "000000";
        when "0001011100010" => rgb <= "100000";
        when "0001011100011" => rgb <= "100000";
        when "0001011100100" => rgb <= "100000";
        when "0001011100101" => rgb <= "100000";
        when "0001011100110" => rgb <= "100000";
        when "0001011100111" => rgb <= "000000";
        when "0001100000000" => rgb <= "000000";
        when "0001100000001" => rgb <= "000000";
        when "0001100000010" => rgb <= "000000";
        when "0001100000011" => rgb <= "000000";
        when "0001100000100" => rgb <= "000000";
        when "0001100000101" => rgb <= "000000";
        when "0001100000110" => rgb <= "000000";
        when "0001100000111" => rgb <= "000000";
        when "0001100001000" => rgb <= "000000";
        when "0001100001001" => rgb <= "000000";
        when "0001100001010" => rgb <= "000000";
        when "0001100001011" => rgb <= "000000";
        when "0001100001100" => rgb <= "000000";
        when "0001100001101" => rgb <= "000000";
        when "0001100001110" => rgb <= "000000";
        when "0001100001111" => rgb <= "000000";
        when "0001100010000" => rgb <= "000000";
        when "0001100010001" => rgb <= "000000";
        when "0001100010010" => rgb <= "000000";
        when "0001100010011" => rgb <= "000000";
        when "0001100010100" => rgb <= "000000";
        when "0001100010101" => rgb <= "000000";
        when "0001100010110" => rgb <= "000000";
        when "0001100010111" => rgb <= "000000";
        when "0001100011000" => rgb <= "000000";
        when "0001100011001" => rgb <= "000000";
        when "0001100011010" => rgb <= "000000";
        when "0001100011011" => rgb <= "000000";
        when "0001100011100" => rgb <= "000000";
        when "0001100011101" => rgb <= "000000";
        when "0001100011110" => rgb <= "000000";
        when "0001100011111" => rgb <= "000000";
        when "0001100100000" => rgb <= "000000";
        when "0001100100001" => rgb <= "000000";
        when "0001100100010" => rgb <= "000000";
        when "0001100100011" => rgb <= "000000";
        when "0001100100100" => rgb <= "000000";
        when "0001100100101" => rgb <= "000000";
        when "0001100100110" => rgb <= "000000";
        when "0001100100111" => rgb <= "000000";
        when "0001101000000" => rgb <= "000000";
        when "0001101000001" => rgb <= "000000";
        when "0001101000010" => rgb <= "000000";
        when "0001101000011" => rgb <= "000000";
        when "0001101000100" => rgb <= "000000";
        when "0001101000101" => rgb <= "000000";
        when "0001101000110" => rgb <= "000000";
        when "0001101000111" => rgb <= "000000";
        when "0001101001000" => rgb <= "000000";
        when "0001101001001" => rgb <= "000000";
        when "0001101001010" => rgb <= "000000";
        when "0001101001011" => rgb <= "000000";
        when "0001101001100" => rgb <= "000000";
        when "0001101001101" => rgb <= "000000";
        when "0001101001110" => rgb <= "000000";
        when "0001101001111" => rgb <= "000000";
        when "0001101010000" => rgb <= "000000";
        when "0001101010001" => rgb <= "000000";
        when "0001101010010" => rgb <= "000000";
        when "0001101010011" => rgb <= "000000";
        when "0001101010100" => rgb <= "000000";
        when "0001101010101" => rgb <= "000000";
        when "0001101010110" => rgb <= "000000";
        when "0001101010111" => rgb <= "000000";
        when "0001101011000" => rgb <= "000000";
        when "0001101011001" => rgb <= "000000";
        when "0001101011010" => rgb <= "000000";
        when "0001101011011" => rgb <= "000000";
        when "0001101011100" => rgb <= "000000";
        when "0001101011101" => rgb <= "000000";
        when "0001101011110" => rgb <= "000000";
        when "0001101011111" => rgb <= "000000";
        when "0001101100000" => rgb <= "000000";
        when "0001101100001" => rgb <= "000000";
        when "0001101100010" => rgb <= "000000";
        when "0001101100011" => rgb <= "000000";
        when "0001101100100" => rgb <= "000000";
        when "0001101100101" => rgb <= "000000";
        when "0001101100110" => rgb <= "000000";
        when "0001101100111" => rgb <= "000000";
        when "0001110000000" => rgb <= "000000";
        when "0001110000001" => rgb <= "000000";
        when "0001110000010" => rgb <= "000000";
        when "0001110000011" => rgb <= "000000";
        when "0001110000100" => rgb <= "000000";
        when "0001110000101" => rgb <= "000000";
        when "0001110000110" => rgb <= "000000";
        when "0001110000111" => rgb <= "000000";
        when "0001110001000" => rgb <= "000000";
        when "0001110001001" => rgb <= "000000";
        when "0001110001010" => rgb <= "000000";
        when "0001110001011" => rgb <= "000000";
        when "0001110001100" => rgb <= "000000";
        when "0001110001101" => rgb <= "000000";
        when "0001110001110" => rgb <= "000000";
        when "0001110001111" => rgb <= "000000";
        when "0001110010000" => rgb <= "000000";
        when "0001110010001" => rgb <= "000000";
        when "0001110010010" => rgb <= "000000";
        when "0001110010011" => rgb <= "000000";
        when "0001110010100" => rgb <= "000000";
        when "0001110010101" => rgb <= "000000";
        when "0001110010110" => rgb <= "000000";
        when "0001110010111" => rgb <= "000000";
        when "0001110011000" => rgb <= "000000";
        when "0001110011001" => rgb <= "000000";
        when "0001110011010" => rgb <= "000000";
        when "0001110011011" => rgb <= "000000";
        when "0001110011100" => rgb <= "000000";
        when "0001110011101" => rgb <= "000000";
        when "0001110011110" => rgb <= "000000";
        when "0001110011111" => rgb <= "000000";
        when "0001110100000" => rgb <= "000000";
        when "0001110100001" => rgb <= "000000";
        when "0001110100010" => rgb <= "000000";
        when "0001110100011" => rgb <= "000000";
        when "0001110100100" => rgb <= "000000";
        when "0001110100101" => rgb <= "000000";
        when "0001110100110" => rgb <= "000000";
        when "0001110100111" => rgb <= "000000";
        when "0001111000000" => rgb <= "000000";
        when "0001111000001" => rgb <= "000000";
        when "0001111000010" => rgb <= "000000";
        when "0001111000011" => rgb <= "000000";
        when "0001111000100" => rgb <= "000000";
        when "0001111000101" => rgb <= "000000";
        when "0001111000110" => rgb <= "000000";
        when "0001111000111" => rgb <= "100000";
        when "0001111001000" => rgb <= "000000";
        when "0001111001001" => rgb <= "000000";
        when "0001111001010" => rgb <= "000000";
        when "0001111001011" => rgb <= "100000";
        when "0001111001100" => rgb <= "000000";
        when "0001111001101" => rgb <= "000000";
        when "0001111001110" => rgb <= "000000";
        when "0001111001111" => rgb <= "100000";
        when "0001111010000" => rgb <= "000000";
        when "0001111010001" => rgb <= "100000";
        when "0001111010010" => rgb <= "100000";
        when "0001111010011" => rgb <= "100000";
        when "0001111010100" => rgb <= "000000";
        when "0001111010101" => rgb <= "100000";
        when "0001111010110" => rgb <= "100000";
        when "0001111010111" => rgb <= "000000";
        when "0001111011000" => rgb <= "000000";
        when "0001111011001" => rgb <= "000000";
        when "0001111011010" => rgb <= "100000";
        when "0001111011011" => rgb <= "000000";
        when "0001111011100" => rgb <= "000000";
        when "0001111011101" => rgb <= "100000";
        when "0001111011110" => rgb <= "100000";
        when "0001111011111" => rgb <= "100000";
        when "0001111100000" => rgb <= "100000";
        when "0001111100001" => rgb <= "000000";
        when "0001111100010" => rgb <= "000000";
        when "0001111100011" => rgb <= "000000";
        when "0001111100100" => rgb <= "000000";
        when "0001111100101" => rgb <= "000000";
        when "0001111100110" => rgb <= "000000";
        when "0001111100111" => rgb <= "000000";
        when "0010000000000" => rgb <= "000000";
        when "0010000000001" => rgb <= "000000";
        when "0010000000010" => rgb <= "000000";
        when "0010000000011" => rgb <= "000000";
        when "0010000000100" => rgb <= "000000";
        when "0010000000101" => rgb <= "000000";
        when "0010000000110" => rgb <= "000000";
        when "0010000000111" => rgb <= "100000";
        when "0010000001000" => rgb <= "000000";
        when "0010000001001" => rgb <= "000000";
        when "0010000001010" => rgb <= "000000";
        when "0010000001011" => rgb <= "100000";
        when "0010000001100" => rgb <= "000000";
        when "0010000001101" => rgb <= "000000";
        when "0010000001110" => rgb <= "000000";
        when "0010000001111" => rgb <= "100000";
        when "0010000010000" => rgb <= "000000";
        when "0010000010001" => rgb <= "000000";
        when "0010000010010" => rgb <= "100000";
        when "0010000010011" => rgb <= "000000";
        when "0010000010100" => rgb <= "000000";
        when "0010000010101" => rgb <= "100000";
        when "0010000010110" => rgb <= "100000";
        when "0010000010111" => rgb <= "000000";
        when "0010000011000" => rgb <= "000000";
        when "0010000011001" => rgb <= "000000";
        when "0010000011010" => rgb <= "100000";
        when "0010000011011" => rgb <= "000000";
        when "0010000011100" => rgb <= "100000";
        when "0010000011101" => rgb <= "000000";
        when "0010000011110" => rgb <= "000000";
        when "0010000011111" => rgb <= "000000";
        when "0010000100000" => rgb <= "000000";
        when "0010000100001" => rgb <= "000000";
        when "0010000100010" => rgb <= "000000";
        when "0010000100011" => rgb <= "000000";
        when "0010000100100" => rgb <= "000000";
        when "0010000100101" => rgb <= "000000";
        when "0010000100110" => rgb <= "000000";
        when "0010000100111" => rgb <= "000000";
        when "0010001000000" => rgb <= "000000";
        when "0010001000001" => rgb <= "000000";
        when "0010001000010" => rgb <= "000000";
        when "0010001000011" => rgb <= "000000";
        when "0010001000100" => rgb <= "000000";
        when "0010001000101" => rgb <= "000000";
        when "0010001000110" => rgb <= "000000";
        when "0010001000111" => rgb <= "100000";
        when "0010001001000" => rgb <= "000000";
        when "0010001001001" => rgb <= "000000";
        when "0010001001010" => rgb <= "000000";
        when "0010001001011" => rgb <= "100000";
        when "0010001001100" => rgb <= "000000";
        when "0010001001101" => rgb <= "000000";
        when "0010001001110" => rgb <= "000000";
        when "0010001001111" => rgb <= "100000";
        when "0010001010000" => rgb <= "000000";
        when "0010001010001" => rgb <= "000000";
        when "0010001010010" => rgb <= "100000";
        when "0010001010011" => rgb <= "000000";
        when "0010001010100" => rgb <= "000000";
        when "0010001010101" => rgb <= "100000";
        when "0010001010110" => rgb <= "000000";
        when "0010001010111" => rgb <= "100000";
        when "0010001011000" => rgb <= "000000";
        when "0010001011001" => rgb <= "000000";
        when "0010001011010" => rgb <= "100000";
        when "0010001011011" => rgb <= "000000";
        when "0010001011100" => rgb <= "100000";
        when "0010001011101" => rgb <= "000000";
        when "0010001011110" => rgb <= "000000";
        when "0010001011111" => rgb <= "000000";
        when "0010001100000" => rgb <= "000000";
        when "0010001100001" => rgb <= "000000";
        when "0010001100010" => rgb <= "000000";
        when "0010001100011" => rgb <= "000000";
        when "0010001100100" => rgb <= "000000";
        when "0010001100101" => rgb <= "000000";
        when "0010001100110" => rgb <= "000000";
        when "0010001100111" => rgb <= "000000";
        when "0010010000000" => rgb <= "000000";
        when "0010010000001" => rgb <= "000000";
        when "0010010000010" => rgb <= "000000";
        when "0010010000011" => rgb <= "000000";
        when "0010010000100" => rgb <= "000000";
        when "0010010000101" => rgb <= "000000";
        when "0010010000110" => rgb <= "000000";
        when "0010010000111" => rgb <= "000000";
        when "0010010001000" => rgb <= "100000";
        when "0010010001001" => rgb <= "000000";
        when "0010010001010" => rgb <= "100000";
        when "0010010001011" => rgb <= "000000";
        when "0010010001100" => rgb <= "100000";
        when "0010010001101" => rgb <= "000000";
        when "0010010001110" => rgb <= "100000";
        when "0010010001111" => rgb <= "000000";
        when "0010010010000" => rgb <= "000000";
        when "0010010010001" => rgb <= "000000";
        when "0010010010010" => rgb <= "100000";
        when "0010010010011" => rgb <= "000000";
        when "0010010010100" => rgb <= "000000";
        when "0010010010101" => rgb <= "100000";
        when "0010010010110" => rgb <= "000000";
        when "0010010010111" => rgb <= "100000";
        when "0010010011000" => rgb <= "000000";
        when "0010010011001" => rgb <= "000000";
        when "0010010011010" => rgb <= "100000";
        when "0010010011011" => rgb <= "000000";
        when "0010010011100" => rgb <= "000000";
        when "0010010011101" => rgb <= "100000";
        when "0010010011110" => rgb <= "100000";
        when "0010010011111" => rgb <= "100000";
        when "0010010100000" => rgb <= "000000";
        when "0010010100001" => rgb <= "000000";
        when "0010010100010" => rgb <= "000000";
        when "0010010100011" => rgb <= "000000";
        when "0010010100100" => rgb <= "000000";
        when "0010010100101" => rgb <= "000000";
        when "0010010100110" => rgb <= "000000";
        when "0010010100111" => rgb <= "000000";
        when "0010011000000" => rgb <= "000000";
        when "0010011000001" => rgb <= "000000";
        when "0010011000010" => rgb <= "000000";
        when "0010011000011" => rgb <= "000000";
        when "0010011000100" => rgb <= "000000";
        when "0010011000101" => rgb <= "000000";
        when "0010011000110" => rgb <= "000000";
        when "0010011000111" => rgb <= "000000";
        when "0010011001000" => rgb <= "100000";
        when "0010011001001" => rgb <= "000000";
        when "0010011001010" => rgb <= "100000";
        when "0010011001011" => rgb <= "000000";
        when "0010011001100" => rgb <= "100000";
        when "0010011001101" => rgb <= "000000";
        when "0010011001110" => rgb <= "100000";
        when "0010011001111" => rgb <= "000000";
        when "0010011010000" => rgb <= "000000";
        when "0010011010001" => rgb <= "000000";
        when "0010011010010" => rgb <= "100000";
        when "0010011010011" => rgb <= "000000";
        when "0010011010100" => rgb <= "000000";
        when "0010011010101" => rgb <= "100000";
        when "0010011010110" => rgb <= "000000";
        when "0010011010111" => rgb <= "000000";
        when "0010011011000" => rgb <= "100000";
        when "0010011011001" => rgb <= "000000";
        when "0010011011010" => rgb <= "100000";
        when "0010011011011" => rgb <= "000000";
        when "0010011011100" => rgb <= "000000";
        when "0010011011101" => rgb <= "000000";
        when "0010011011110" => rgb <= "000000";
        when "0010011011111" => rgb <= "000000";
        when "0010011100000" => rgb <= "100000";
        when "0010011100001" => rgb <= "000000";
        when "0010011100010" => rgb <= "000000";
        when "0010011100011" => rgb <= "000000";
        when "0010011100100" => rgb <= "000000";
        when "0010011100101" => rgb <= "000000";
        when "0010011100110" => rgb <= "000000";
        when "0010011100111" => rgb <= "000000";
        when "0010100000000" => rgb <= "000000";
        when "0010100000001" => rgb <= "000000";
        when "0010100000010" => rgb <= "000000";
        when "0010100000011" => rgb <= "000000";
        when "0010100000100" => rgb <= "000000";
        when "0010100000101" => rgb <= "000000";
        when "0010100000110" => rgb <= "000000";
        when "0010100000111" => rgb <= "000000";
        when "0010100001000" => rgb <= "100000";
        when "0010100001001" => rgb <= "000000";
        when "0010100001010" => rgb <= "100000";
        when "0010100001011" => rgb <= "000000";
        when "0010100001100" => rgb <= "100000";
        when "0010100001101" => rgb <= "000000";
        when "0010100001110" => rgb <= "100000";
        when "0010100001111" => rgb <= "000000";
        when "0010100010000" => rgb <= "000000";
        when "0010100010001" => rgb <= "000000";
        when "0010100010010" => rgb <= "100000";
        when "0010100010011" => rgb <= "000000";
        when "0010100010100" => rgb <= "000000";
        when "0010100010101" => rgb <= "100000";
        when "0010100010110" => rgb <= "000000";
        when "0010100010111" => rgb <= "000000";
        when "0010100011000" => rgb <= "100000";
        when "0010100011001" => rgb <= "000000";
        when "0010100011010" => rgb <= "100000";
        when "0010100011011" => rgb <= "000000";
        when "0010100011100" => rgb <= "000000";
        when "0010100011101" => rgb <= "000000";
        when "0010100011110" => rgb <= "000000";
        when "0010100011111" => rgb <= "000000";
        when "0010100100000" => rgb <= "100000";
        when "0010100100001" => rgb <= "000000";
        when "0010100100010" => rgb <= "000000";
        when "0010100100011" => rgb <= "000000";
        when "0010100100100" => rgb <= "000000";
        when "0010100100101" => rgb <= "000000";
        when "0010100100110" => rgb <= "000000";
        when "0010100100111" => rgb <= "000000";
        when "0010101000000" => rgb <= "000000";
        when "0010101000001" => rgb <= "000000";
        when "0010101000010" => rgb <= "000000";
        when "0010101000011" => rgb <= "000000";
        when "0010101000100" => rgb <= "000000";
        when "0010101000101" => rgb <= "000000";
        when "0010101000110" => rgb <= "000000";
        when "0010101000111" => rgb <= "000000";
        when "0010101001000" => rgb <= "000000";
        when "0010101001001" => rgb <= "100000";
        when "0010101001010" => rgb <= "000000";
        when "0010101001011" => rgb <= "000000";
        when "0010101001100" => rgb <= "000000";
        when "0010101001101" => rgb <= "100000";
        when "0010101001110" => rgb <= "000000";
        when "0010101001111" => rgb <= "000000";
        when "0010101010000" => rgb <= "000000";
        when "0010101010001" => rgb <= "000000";
        when "0010101010010" => rgb <= "100000";
        when "0010101010011" => rgb <= "000000";
        when "0010101010100" => rgb <= "000000";
        when "0010101010101" => rgb <= "100000";
        when "0010101010110" => rgb <= "000000";
        when "0010101010111" => rgb <= "000000";
        when "0010101011000" => rgb <= "000000";
        when "0010101011001" => rgb <= "100000";
        when "0010101011010" => rgb <= "100000";
        when "0010101011011" => rgb <= "000000";
        when "0010101011100" => rgb <= "000000";
        when "0010101011101" => rgb <= "000000";
        when "0010101011110" => rgb <= "000000";
        when "0010101011111" => rgb <= "000000";
        when "0010101100000" => rgb <= "100000";
        when "0010101100001" => rgb <= "000000";
        when "0010101100010" => rgb <= "000000";
        when "0010101100011" => rgb <= "000000";
        when "0010101100100" => rgb <= "000000";
        when "0010101100101" => rgb <= "000000";
        when "0010101100110" => rgb <= "000000";
        when "0010101100111" => rgb <= "000000";
        when "0010110000000" => rgb <= "000000";
        when "0010110000001" => rgb <= "000000";
        when "0010110000010" => rgb <= "000000";
        when "0010110000011" => rgb <= "000000";
        when "0010110000100" => rgb <= "000000";
        when "0010110000101" => rgb <= "000000";
        when "0010110000110" => rgb <= "000000";
        when "0010110000111" => rgb <= "000000";
        when "0010110001000" => rgb <= "000000";
        when "0010110001001" => rgb <= "100000";
        when "0010110001010" => rgb <= "000000";
        when "0010110001011" => rgb <= "000000";
        when "0010110001100" => rgb <= "000000";
        when "0010110001101" => rgb <= "100000";
        when "0010110001110" => rgb <= "000000";
        when "0010110001111" => rgb <= "000000";
        when "0010110010000" => rgb <= "000000";
        when "0010110010001" => rgb <= "100000";
        when "0010110010010" => rgb <= "100000";
        when "0010110010011" => rgb <= "100000";
        when "0010110010100" => rgb <= "000000";
        when "0010110010101" => rgb <= "100000";
        when "0010110010110" => rgb <= "000000";
        when "0010110010111" => rgb <= "000000";
        when "0010110011000" => rgb <= "000000";
        when "0010110011001" => rgb <= "100000";
        when "0010110011010" => rgb <= "100000";
        when "0010110011011" => rgb <= "000000";
        when "0010110011100" => rgb <= "100000";
        when "0010110011101" => rgb <= "100000";
        when "0010110011110" => rgb <= "100000";
        when "0010110011111" => rgb <= "100000";
        when "0010110100000" => rgb <= "000000";
        when "0010110100001" => rgb <= "000000";
        when "0010110100010" => rgb <= "000000";
        when "0010110100011" => rgb <= "000000";
        when "0010110100100" => rgb <= "000000";
        when "0010110100101" => rgb <= "000000";
        when "0010110100110" => rgb <= "000000";
        when "0010110100111" => rgb <= "000000";
        when "0010111000000" => rgb <= "000000";
        when "0010111000001" => rgb <= "000000";
        when "0010111000010" => rgb <= "000000";
        when "0010111000011" => rgb <= "000000";
        when "0010111000100" => rgb <= "000000";
        when "0010111000101" => rgb <= "000000";
        when "0010111000110" => rgb <= "000000";
        when "0010111000111" => rgb <= "000000";
        when "0010111001000" => rgb <= "000000";
        when "0010111001001" => rgb <= "000000";
        when "0010111001010" => rgb <= "000000";
        when "0010111001011" => rgb <= "000000";
        when "0010111001100" => rgb <= "000000";
        when "0010111001101" => rgb <= "000000";
        when "0010111001110" => rgb <= "000000";
        when "0010111001111" => rgb <= "000000";
        when "0010111010000" => rgb <= "000000";
        when "0010111010001" => rgb <= "000000";
        when "0010111010010" => rgb <= "000000";
        when "0010111010011" => rgb <= "000000";
        when "0010111010100" => rgb <= "000000";
        when "0010111010101" => rgb <= "000000";
        when "0010111010110" => rgb <= "000000";
        when "0010111010111" => rgb <= "000000";
        when "0010111011000" => rgb <= "000000";
        when "0010111011001" => rgb <= "000000";
        when "0010111011010" => rgb <= "000000";
        when "0010111011011" => rgb <= "000000";
        when "0010111011100" => rgb <= "000000";
        when "0010111011101" => rgb <= "000000";
        when "0010111011110" => rgb <= "000000";
        when "0010111011111" => rgb <= "000000";
        when "0010111100000" => rgb <= "000000";
        when "0010111100001" => rgb <= "000000";
        when "0010111100010" => rgb <= "000000";
        when "0010111100011" => rgb <= "000000";
        when "0010111100100" => rgb <= "000000";
        when "0010111100101" => rgb <= "000000";
        when "0010111100110" => rgb <= "000000";
        when "0010111100111" => rgb <= "000000";
        when "0011000000000" => rgb <= "000000";
        when "0011000000001" => rgb <= "000000";
        when "0011000000010" => rgb <= "000000";
        when "0011000000011" => rgb <= "000000";
        when "0011000000100" => rgb <= "000000";
        when "0011000000101" => rgb <= "000000";
        when "0011000000110" => rgb <= "000000";
        when "0011000000111" => rgb <= "000000";
        when "0011000001000" => rgb <= "000000";
        when "0011000001001" => rgb <= "000000";
        when "0011000001010" => rgb <= "000000";
        when "0011000001011" => rgb <= "000000";
        when "0011000001100" => rgb <= "000000";
        when "0011000001101" => rgb <= "000000";
        when "0011000001110" => rgb <= "000000";
        when "0011000001111" => rgb <= "000000";
        when "0011000010000" => rgb <= "000000";
        when "0011000010001" => rgb <= "000000";
        when "0011000010010" => rgb <= "000000";
        when "0011000010011" => rgb <= "000000";
        when "0011000010100" => rgb <= "000000";
        when "0011000010101" => rgb <= "000000";
        when "0011000010110" => rgb <= "000000";
        when "0011000010111" => rgb <= "000000";
        when "0011000011000" => rgb <= "000000";
        when "0011000011001" => rgb <= "000000";
        when "0011000011010" => rgb <= "000000";
        when "0011000011011" => rgb <= "000000";
        when "0011000011100" => rgb <= "000000";
        when "0011000011101" => rgb <= "000000";
        when "0011000011110" => rgb <= "000000";
        when "0011000011111" => rgb <= "000000";
        when "0011000100000" => rgb <= "000000";
        when "0011000100001" => rgb <= "000000";
        when "0011000100010" => rgb <= "000000";
        when "0011000100011" => rgb <= "000000";
        when "0011000100100" => rgb <= "000000";
        when "0011000100101" => rgb <= "000000";
        when "0011000100110" => rgb <= "000000";
        when "0011000100111" => rgb <= "000000";
        when "0011001000000" => rgb <= "000000";
        when "0011001000001" => rgb <= "000000";
        when "0011001000010" => rgb <= "000000";
        when "0011001000011" => rgb <= "000000";
        when "0011001000100" => rgb <= "000000";
        when "0011001000101" => rgb <= "000000";
        when "0011001000110" => rgb <= "000000";
        when "0011001000111" => rgb <= "000000";
        when "0011001001000" => rgb <= "000000";
        when "0011001001001" => rgb <= "000000";
        when "0011001001010" => rgb <= "000000";
        when "0011001001011" => rgb <= "000000";
        when "0011001001100" => rgb <= "000000";
        when "0011001001101" => rgb <= "000000";
        when "0011001001110" => rgb <= "000000";
        when "0011001001111" => rgb <= "000000";
        when "0011001010000" => rgb <= "000000";
        when "0011001010001" => rgb <= "000000";
        when "0011001010010" => rgb <= "000000";
        when "0011001010011" => rgb <= "000000";
        when "0011001010100" => rgb <= "000000";
        when "0011001010101" => rgb <= "000000";
        when "0011001010110" => rgb <= "000000";
        when "0011001010111" => rgb <= "000000";
        when "0011001011000" => rgb <= "000000";
        when "0011001011001" => rgb <= "000000";
        when "0011001011010" => rgb <= "000000";
        when "0011001011011" => rgb <= "000000";
        when "0011001011100" => rgb <= "000000";
        when "0011001011101" => rgb <= "000000";
        when "0011001011110" => rgb <= "000000";
        when "0011001011111" => rgb <= "000000";
        when "0011001100000" => rgb <= "000000";
        when "0011001100001" => rgb <= "000000";
        when "0011001100010" => rgb <= "000000";
        when "0011001100011" => rgb <= "000000";
        when "0011001100100" => rgb <= "000000";
        when "0011001100101" => rgb <= "000000";
        when "0011001100110" => rgb <= "000000";
        when "0011001100111" => rgb <= "000000";
        when "0011010000000" => rgb <= "000000";
        when "0011010000001" => rgb <= "000000";
        when "0011010000010" => rgb <= "000000";
        when "0011010000011" => rgb <= "000000";
        when "0011010000100" => rgb <= "000000";
        when "0011010000101" => rgb <= "000000";
        when "0011010000110" => rgb <= "000000";
        when "0011010000111" => rgb <= "000000";
        when "0011010001000" => rgb <= "000000";
        when "0011010001001" => rgb <= "000000";
        when "0011010001010" => rgb <= "000000";
        when "0011010001011" => rgb <= "000000";
        when "0011010001100" => rgb <= "000000";
        when "0011010001101" => rgb <= "000000";
        when "0011010001110" => rgb <= "000000";
        when "0011010001111" => rgb <= "000000";
        when "0011010010000" => rgb <= "000000";
        when "0011010010001" => rgb <= "000000";
        when "0011010010010" => rgb <= "000000";
        when "0011010010011" => rgb <= "000000";
        when "0011010010100" => rgb <= "000000";
        when "0011010010101" => rgb <= "000000";
        when "0011010010110" => rgb <= "000000";
        when "0011010010111" => rgb <= "000000";
        when "0011010011000" => rgb <= "000000";
        when "0011010011001" => rgb <= "000000";
        when "0011010011010" => rgb <= "000000";
        when "0011010011011" => rgb <= "000000";
        when "0011010011100" => rgb <= "000000";
        when "0011010011101" => rgb <= "000000";
        when "0011010011110" => rgb <= "000000";
        when "0011010011111" => rgb <= "000000";
        when "0011010100000" => rgb <= "000000";
        when "0011010100001" => rgb <= "000000";
        when "0011010100010" => rgb <= "000000";
        when "0011010100011" => rgb <= "000000";
        when "0011010100100" => rgb <= "000000";
        when "0011010100101" => rgb <= "000000";
        when "0011010100110" => rgb <= "000000";
        when "0011010100111" => rgb <= "000000";
        when "0011011000000" => rgb <= "000000";
        when "0011011000001" => rgb <= "000000";
        when "0011011000010" => rgb <= "000000";
        when "0011011000011" => rgb <= "000000";
        when "0011011000100" => rgb <= "000000";
        when "0011011000101" => rgb <= "000000";
        when "0011011000110" => rgb <= "000000";
        when "0011011000111" => rgb <= "000000";
        when "0011011001000" => rgb <= "000000";
        when "0011011001001" => rgb <= "000000";
        when "0011011001010" => rgb <= "000000";
        when "0011011001011" => rgb <= "000000";
        when "0011011001100" => rgb <= "000000";
        when "0011011001101" => rgb <= "000000";
        when "0011011001110" => rgb <= "000000";
        when "0011011001111" => rgb <= "000000";
        when "0011011010000" => rgb <= "000000";
        when "0011011010001" => rgb <= "000000";
        when "0011011010010" => rgb <= "000000";
        when "0011011010011" => rgb <= "000000";
        when "0011011010100" => rgb <= "000000";
        when "0011011010101" => rgb <= "000000";
        when "0011011010110" => rgb <= "000000";
        when "0011011010111" => rgb <= "000000";
        when "0011011011000" => rgb <= "000000";
        when "0011011011001" => rgb <= "000000";
        when "0011011011010" => rgb <= "000000";
        when "0011011011011" => rgb <= "000000";
        when "0011011011100" => rgb <= "000000";
        when "0011011011101" => rgb <= "000000";
        when "0011011011110" => rgb <= "000000";
        when "0011011011111" => rgb <= "000000";
        when "0011011100000" => rgb <= "000000";
        when "0011011100001" => rgb <= "000000";
        when "0011011100010" => rgb <= "000000";
        when "0011011100011" => rgb <= "000000";
        when "0011011100100" => rgb <= "000000";
        when "0011011100101" => rgb <= "000000";
        when "0011011100110" => rgb <= "000000";
        when "0011011100111" => rgb <= "000000";
        when "0011100000000" => rgb <= "000000";
        when "0011100000001" => rgb <= "000000";
        when "0011100000010" => rgb <= "000000";
        when "0011100000011" => rgb <= "000000";
        when "0011100000100" => rgb <= "000000";
        when "0011100000101" => rgb <= "000000";
        when "0011100000110" => rgb <= "000000";
        when "0011100000111" => rgb <= "000000";
        when "0011100001000" => rgb <= "000000";
        when "0011100001001" => rgb <= "000000";
        when "0011100001010" => rgb <= "000000";
        when "0011100001011" => rgb <= "000000";
        when "0011100001100" => rgb <= "000000";
        when "0011100001101" => rgb <= "000000";
        when "0011100001110" => rgb <= "000000";
        when "0011100001111" => rgb <= "000000";
        when "0011100010000" => rgb <= "000000";
        when "0011100010001" => rgb <= "000000";
        when "0011100010010" => rgb <= "000000";
        when "0011100010011" => rgb <= "000000";
        when "0011100010100" => rgb <= "000000";
        when "0011100010101" => rgb <= "000000";
        when "0011100010110" => rgb <= "000000";
        when "0011100010111" => rgb <= "000000";
        when "0011100011000" => rgb <= "000000";
        when "0011100011001" => rgb <= "000000";
        when "0011100011010" => rgb <= "000000";
        when "0011100011011" => rgb <= "000000";
        when "0011100011100" => rgb <= "000000";
        when "0011100011101" => rgb <= "000000";
        when "0011100011110" => rgb <= "000000";
        when "0011100011111" => rgb <= "000000";
        when "0011100100000" => rgb <= "000000";
        when "0011100100001" => rgb <= "000000";
        when "0011100100010" => rgb <= "000000";
        when "0011100100011" => rgb <= "000000";
        when "0011100100100" => rgb <= "000000";
        when "0011100100101" => rgb <= "000000";
        when "0011100100110" => rgb <= "000000";
        when "0011100100111" => rgb <= "000000";
        when "0011101000000" => rgb <= "000000";
        when "0011101000001" => rgb <= "000000";
        when "0011101000010" => rgb <= "000000";
        when "0011101000011" => rgb <= "000000";
        when "0011101000100" => rgb <= "000000";
        when "0011101000101" => rgb <= "000000";
        when "0011101000110" => rgb <= "000000";
        when "0011101000111" => rgb <= "000000";
        when "0011101001000" => rgb <= "000000";
        when "0011101001001" => rgb <= "000000";
        when "0011101001010" => rgb <= "000000";
        when "0011101001011" => rgb <= "000000";
        when "0011101001100" => rgb <= "000000";
        when "0011101001101" => rgb <= "000000";
        when "0011101001110" => rgb <= "000000";
        when "0011101001111" => rgb <= "000000";
        when "0011101010000" => rgb <= "000000";
        when "0011101010001" => rgb <= "000000";
        when "0011101010010" => rgb <= "000000";
        when "0011101010011" => rgb <= "000000";
        when "0011101010100" => rgb <= "000000";
        when "0011101010101" => rgb <= "000000";
        when "0011101010110" => rgb <= "000000";
        when "0011101010111" => rgb <= "000000";
        when "0011101011000" => rgb <= "000000";
        when "0011101011001" => rgb <= "000000";
        when "0011101011010" => rgb <= "000000";
        when "0011101011011" => rgb <= "000000";
        when "0011101011100" => rgb <= "000000";
        when "0011101011101" => rgb <= "000000";
        when "0011101011110" => rgb <= "000000";
        when "0011101011111" => rgb <= "000000";
        when "0011101100000" => rgb <= "000000";
        when "0011101100001" => rgb <= "000000";
        when "0011101100010" => rgb <= "000000";
        when "0011101100011" => rgb <= "000000";
        when "0011101100100" => rgb <= "000000";
        when "0011101100101" => rgb <= "000000";
        when "0011101100110" => rgb <= "000000";
        when "0011101100111" => rgb <= "000000";
        when others => rgb <= "000000";
            end case;
end if;
	end process;
	   totaladr <= std_logic_vector(y_cord) & std_logic_vector(x_cord);
end;